��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X������r��#@�/�����4�p5���4;Od��N��r�I#��7h��$�(��?�g:�ZGY�bӍ��0Yzb0o �Β��A���p�6� �����4���e����7�5G��Ξ@��/6����=;+�Cgt�ܫ����ߥo��yqa�ĝ!�G�F#{5� �E؃��\il����A�E�sƸ��]��i��Y���i���	��'i�6�9U�x� ��n���}FA3>[4��L�������g�l�Ju�;�I~m_��dA�e$�)�R��SI�m����[&�wY��m��5�qKhFZ\ϵ�+��	%lke��%�Y�C_V��Y��
tzP���ܫ�FR�34������a_���[B솋���UX��\��t��ň@�%>&��YүLIH<%��/E�5x��v��/&�#X#/��u��Jf�Hh���Q�8�=[����������γA�Ni�0?ut�"�/{.�g��?FڟBڳ�w��� ?����P��Ø������$�GN&>�~g�"���.���V@i�9M���D�::�l�����u�gy&���ROF�� `{�B�YD�,$�^���w���oHH���{}��/�<ŗ����Z�F�~�:��i)�|�W�B��c�C֏�v�����8-4UP��3�0���=�5ި$�T���?�"� ��+��o6��fG�a]_�Lw�Sa�iN�x[�ǔ�ظ8���ʐ@j���Zf�Tt�cv���OM0�ƥ�>C� x;��P&@��Y�&9jI%d�Zk�-�h�K&�����u]��Ln�]�-��5�u^~����j*T�~N�Wv�>�i�8�a�d��`�qVL��Ok����=8�T�<�(�����T�<�"8.U�AOW���e�����%6��"�Ij�S�{o*���
$+�f]n�]�.ǀO��~�х����y�~���	D&crQv���� Fi��-�ƒGcJ
���@�A��ëjВP��X��@���ٶ#��@���Eq��M�\��Ÿ`�`zr��5RK�����tk �#)��Aq�r�Sg#����oֹe�8�S�U��k���=��V5� �A�=��� 4;\��I��z��	��%9F�zmV�+��5�8ܫ��ҷD�plc��,���L�����B�����J�b����x��3a0��N�V���(4H�ʼ�_��?��.�f�J�~���I�<j�|a�9Q�a��}�����	��,~H۪Q����gⅠ�~�����B��	����:$��p�σ���f�ҫ��z���oS��Ԭ��z#U��@�>��x���rX�M�u2��cs1���)��yO8*�SdX
��еI"k+My+����/� O�|E̯$���X����?�̓q�V�Jxe�����
6�F!�Єh0����<��"��[Ne�⍮�y}��[��ن���s,�%�
�k$�&��V���k6mp���+d���b�Q�IQ�r�	{Q��ݞ�l}���&�כ���v:냉�3�o��m�-�e��k��!��A��b��?~�-�j:���LD~��0�y+@�մ�Q�R��{7�l��WH[�
$(�SA����!Q~�#z����q�:�jj˴K�n��|*|_�+�5���o����&�F�eٵڜw�8/�U�L��XW��I���_���ol��uR�F��)ï����q��V6�5l�~���]����o�p�RuXb��κ�;�g������w�>�ɫ����r�D�el ��"*� �W���=&�e���!2�@XS��a@Z2)�{�^�q!���F�p��^��?!�>A�^�qH��H�̚��{{��J�ϡж�.�)~6-q� ��� � �J��Ѳ+�~��S��Fgo�p#�ώ����@�����F�]��$��w�,5Y�"��'�̃�+��� ����1_'�P�PG�l�ׂ	O#4��4�[O�?���\�k?����|a��"���_���C�bY�.k��L�Vy�M�`��?������h�V��v0|�<.C���	O�	��B�RV9�(��[�y�"dp�0]#HֱYP�j��nX_cd�Kj|,�1cD�>hC�Ŝ}��9��}l]�n�m�����G�J.%]�wa��"�m\�\@�S�T�V�o�z��Ga,Xl���٘��K9d�(�V�E�iIx� m�m?���jy��0����bl`����ܼ���`'$��J-:���O�TಀF�]��AP�ϥ�@F��;Mbu��5�~��Ko�|&��
�@R@`���I��eEo�ɶ��p�M�	 o���.�]�?s��uuu%��� ���u��ѾJ}Ar�l0�3H�W��e�����ce���3 �V�Kã���z�(�VY�.�$��������vq����hR�@8���N��?���#7q|Rn!��-(Э�d�PZD���#N�
�lkn�cr��(1��&6ВКr.�:B?·�8>3�f�L�ˍ�@�9~�X��ȯ?xa���{%�4��m<q<�������Xf��Ve��� �L��d��R��4:�>e �Vu?�7ӫ�__b21�(��V�o�k���J����h-�� 1qa�<bҥ����{�iw�W���2�,B 2-Uΐ����β"�8���P���P�ʨa�`7��﷭�`�vj��.�{��]�B'o��@�~�$��l��1n��IR���[m�G.��:�e���L��xj
9�FA�)�=�\����� �3��=�a�f�P��
��jm�Ş�Y��Fɾp��`�~;��͗Ȧ�QE;����'fݕ3��x����������"Y2�B�x7���D+�����64f�=�`&��{���u�}��~%s�\8��/�`�Wkq�^r�a4�r=�Ao���%�]!dM�Y'2�N2H��ǻ��V'��������j%�2��ы�0{c�XDfm�����@5��a�-.{μ�]�ya�7���U�.J��	X~����	%pI'�z(h��(�ʲ.����@}�װ4��sV	��Y��ˍ��d��B����!��#9gqh�"'w!���rl�@2?8�������2��t��HIz��yu��S�H��g���:Ɗ�����7k\�c����y1��!�L�-�rٟ��\>5*3��=O#���������*���'��>�4�L��!u�R��awVw�-M�_�1����j�$3I����*�P�C�MC��.����������\�<�H�E�E�u`�	��A�1�������Կ�t�mI5h��\� �����9���g�C����D�W+��o�y-�d�X��h��˚v7BB
�c"�xkT�=��@������^�6�"U�1 �/���(8A�;B�"9Eb�����J44z7����}4���;ت��P켁)f�ZU&4Z��e�Ys{2���6L����<�wf�R�!U���������F߃���Œ��²�h��3��G�幅�f;�<5]/Z��j��Ŏ�>#��Cr�}���O��B�@� �V߶�*J����+���a~5i`�-ھ����4�o���=�q#�#���q]:��zއHba��H;|Z��p"�U�yl�:�a@�K�W�[0�ḓR�ڈ��s��LR>�
�%n��)���F5�s�Ҩ!$4� f���~�;�n�<��l�����hZǸ%��,��C�[_-�3���E���W'���P���A�?��c֡��������H�/��T�_$����R5D�.�n�V*u<��qP��Qn� �Y�&�f� ES>Kּ����޼��MY��Z���NZ ��n1o�A�TNk���b@����Vw�4unN�ܰ�4��Г��=Kp/�5�0ȿv B�s)���� P@�H�c�Pf}j��X�F���(�jRX֘N��D��������^Qp��7�E&��[n|7zʅQ��堚!���9�ōoQto�	FG�,"g�z�n��.��O":-a��";�Q8�h.~u����gsB�����1��Y��Λ�f��7�[L�7���ˑ���|zj�紬YUe�t�E.��R�#���0��.�����	�A�����!g��� TY}�84`иe?�ꤓ�s�j�a���w�("�#�O�b�M��]��8����R�/���I���5�5d����JZ��k�~3��ݸW����8_�l⟙��&HV��+��wk��o�]0���w�����@l�S��.'3ש����`��Dv;	~��I����(��N|�C	��|g ��×���S�Bc58�"����
�<��H\���FRg �S4�rt�W�l��Q�׺��<D�~��������~�8`�v&�jL�w`�贍Q|U�$�Cp�U5uK?��w�^o�� ��R��tq���+�7�P��������
��� n���[z��e�kqZ�va��X�l�7ws�Ѭ)$����
��v�-7�� 6��s0��:�J���6_�R����H�s�q��*4�j*�x�q4P,����*4Z�Ч������4,nb[�<1���z>>�k�>p��%$o��=9�b񺆲i�[�nD"+!�&�7O�f�J���uJ�q3���l[�Z�bz���Yy���o�j�*��O(��4q]A��P>$ǽ7�����)d�e�wt�)������F��m�Gj+,"8���;�?���;ۇ�
�0�Q;w��j`8g���X�d�X�B�.�vC�Y�0�V+
�=BC���`���W����yĭ�N!��!�=�4S/�oo�����
.�g?�r������ޭ��!||��j�_5�ɍ)m!���@�ð���7%��O����M��ץi�]_�x־;ZS?c�tz	���L��؄o�>�$?�WY�5�q����k���5�7�y�" �����l4a��+Z�ts?y��%8%�Ζ��Ta�u�`��[��5W�Ё~�o]��^Q������p�wm�����ei_��r_�VDf,*��s�V��,}#��T����"y��`$X���ک~v(���@�ɋ<�B���l� )�f���$�Q}�Gǰ�u�(�t���o:���0��x��/j�I��M�h�0��w�M��z���0B�I��K��3�mi�-�� ��_���;� �3�A��r��.��+S�$���_&烢��(շ�E�Iqʺ���B}���
K�6c'��7�%�&��1��8h�]puϦ��r� 	"8�M�>��n�΁��k�MYm@�81�ї�I���O	�'��u#=��ߏ[:^5h��ŪU��[�}��B%$V�<������G ����[m�;R��%4���kƊ�y7��u@�୯���4����i��7$��J��E~oG0H�c{2f���ڿ�}K��T�pV8��W�h�(���
���A��QA$r�Cl��
�D�wT{^�E#)���E� �̒%�?V����|�_9���(9�'�G-��R,���G�!�i���6v��� S�VҮ����MG�V�/������S<�g��������|���gXU�0�}�b�`�e��5�K���v}���
����ߣ/�c��8����U/�|��[���G�7��wDչ�L�~��8rf�e���Y%x�Wǲ-.��>b�������4�=mU��5]�����q34�}�vp����|�B�i�C�s�p���@��ºoŃ'����2��[ڂ���:��ki�[�,�s  |s��dW�_��?Jzu�xӨ���YFgn�FR8���K�&{�d�J*ҹ�6�˴�#6߾�sM����yZ�A�V��Ҋ��.!�����x��� �f�"�زD:O�-k3�u-���p�!9j�k\�ϲ��ܝ����È�žpG���zR\�1�(}J˛@ S��Lt���������?�¿��)��)�;#{<+�3���l�dS�T霑��?�t#�StW� h<��Y���&g��n��n�<�1���!zU2ܸ�2�i���7IA����њ��h��
�B^ʨeh�'(�{r6����\f��u�*�!'���^���<D��QS���JPJ��Q7�UVR].�~�*�'�qٖ.R�j��9�5�p��l�n�'Z���Y?9��D&��r�G]s�7�gFbyvJ������T�l�iڝ�L���̬<cs����a�g�sօ�A/mL�Ex��C�0+ �aN���IL����ݵ9�����եﲟ����>*��Q��s�c�j.���I���_��
ُ��o@�R�B]M��!��mY���-V��� }25���`��V^r���1�!'S
��������i
�Ŝ�:Z�� ��;�J'�V2�<���n��rx@�Q�y��K����y\�ǌ-��`��]��.�uO�6D�>�*:�y����a �2�.Q�e��OW/*�����>�V��K0�� ���1��rV�D5���
-H�@<�1��ٍ�gd�:kDx�33�#ރ��E�!�5bG�g�@�>�d���T���A�J�(�m5�ڶͩ��
F�c�8�>Tg��Ft��%�R��"�b���z�s��"m��~���ݙ�@�����<���og�T�J�J!{efeQ7VK��޶V:ɰ ����
��g�$����!�$�pх�e�R�3���cYٺb��k�͏���c��o���]2j�.����+鳚����8Cs%T'�����B���]�Rt�w�x�	�u���^s�c��g�皔*�E^�ֻ�1�<�A(��՝����Hhr��a^�[�_��J�0n��0v^��������<{����+����*:���rvbcKDs�1J��������W�v���x�ﵧ>�:�x�vP��_c�j�/��*]u�WA@v��,#��p���6����8@N���3-21t�����d?'�U�c�����`uoТ�a�w]xlfS:��1�"H�"��=��;*8/+ʠ\���X�A�.GGW@�O+�A:���B�x�������T�it���q��+���L �I1\O�>d�y\H��Z(�X�D�DYMG���a����I�b��;ˍz��C����� +T{��$�L�zl��IMƈ��H�g�ʅ����	=?��JB����1�>]0�$�r?ccAV�W�FG�W����Vc���88�ŏ��kI�(^����B���w�@v܉��ks�⪊]-�|k��W9�1V�J�t��V9�Y�/俁Zs�b��R��;�3j4��DEЙÏV)�Ȼ}�D����Ĵ�1�GG͙�J�[t����e&I��O���h=���]�"1o�\Ԉ�6�ir������]y�XSz����@K�]^ �P!n��2j�����#�L���i�tK�w�{`:c|9���w'�Jo9z�>�*�;~|&P����J�Q�д!�d9AB���e�����ӳ���A�������H�=�B` ��?��w)�ď>>����9���\�;��GPn�$�c$h��]�4�$�&���%��~��m�c*�`��~#(�q��� �����,c�J_��tl7=�W�@�rkb@��p;+���r%��4n4~�6�\�$E'��Wx��h�x��_�G�	.D V���-��q<��_OL��s�t	�=��Tq2#��Bb���?��HL�lb�'dz�Jz�{��](|�ER,��}d�0=�j��)��Iil�U��q6),,䶢?������?�^��*�]tL�pdԌHP��i�_��$�	��g�D�]�6|�E��F�<c!h	�Fi��,�^U��,�	G�@����z]�xj?i"BE�{\�`95yZ����!ݶ�f��a1�u��ȔP�M��i������'�$�ڛ���}uxG��ɇ�IoO�t�ZkM4"Ǎ�QD��j���Q�k��[d��q����M��M���uS`E ƱZg4����[_�UQe�p�J�r��8]`��Q�޿F�V����md|��Q��؜� 0h:.��T�9k-yVY�K�u��T�j4�5\D�`|�E�ɕ�X�~�ܮ�_UK}�F��`��?�+�qTnH�Ot�J.�J`�E�n�<VU;o�Z�6R �A��=��\/X�3	_���`�0~�6TSq����Vɇ�2�&��%!J��6��=���C�����k���vj/7��J9 `�[�N�V��^F���'��-�a�a�%	d����/�VK����uKW5g��4$fJ��T���-԰�j0o΄�@�cpЭpq�
��v�]�#DH5>.сv(����:lq>�J�|� � �����u�3L'���6��>/?��q���'�m������N��aH?Z�����R��H$U��Ј�/���^3���������x��|i�ޯn�ա�(�#�Π�'&��S>O�x�z�5����8��ydE1����:B���3��b�4�z��	����/c���C�m=�w�����B�S(�� <��?����B�(ܭ�7�1�*�4��=k����|g�D��L���,�E%C�R��Ȑeɵ�u�S�Ljoǩ�F�#x�g�XQ�芼':���雘����~�50��XC�gJ�]���;�{�ʚ1�F�i��B�!L`��4��b�C�s4	�
 w	�����qi���[J��3�I�J���cS��\Q��qL��TYEW�A�2��Y����2��S*f����y�����h��΄�S�f����C%\�D�hc��D{��l�P<(�2U�N��_\�ڮ9�;�yP7��!�7t����n8�U�3�W� ��0kR�)�	��UH�P��ũ�r��ٔ�	D@A>��1������>��1.�ݣ/���nb�d���SA_�3�!i�?���-�?l�d�؁~J�Q�-����@�h����&�I��z�:�	�6с��W$J����Z����M[E�FC(��KU�Ib��\+��?���8	k��K@E�A�5׍ fڡ%G~�J��3zF��s�w2	��'�J�v��}��{�`��<���^A�����6>���=�=�a<� �q=E�2 e�ƻ/�X��)���OUs��ݬ��Yf�HA���g}�w8�ȫ8��"�m#���)!# 5�'8�>Կ����ISc��F�%X����Fjc�	J�y̈́��l���C4�͖��@������GRM �	��|T�3|�>����Q��69�zg$�����GÈ��<��+��B��[�G;�>t}xT�='����{�)��{⣱�U �R6�Vs�*i��Qn�xsf��?YA�>�����X���&��������;�,�z�
�be�����s�z~Dm.��qT�F��Ƥ��cyWv3�*��W�}�-ʰte��A��v`�kZv��X���/sꦻ1r�c��uD|���?�^�� �I��+�p�����u�,��0L�eqЗBi������<�M>��_�mm�	�*Q�l}k��\�*S���Ό���b�N��e��s�s���9:r�|��A��s���r��`r�C4�u�ԓ�4��n���S<���Y�9�5�5:�Έ�_���lK�x>�_�a6�T��0��^>O�솥g~�CY\,���%gn$D�t��^
�xVĩF����:��-���lY"-5���jݳ%E��;�}.�w�/Ğ.��m��'���8�|	P΁ �s�f� d2r�=?mi8��6	Y*Z֘j�{ a��Y#�3H��=&��d�V���	G��^#>q/)�ʵwb���~�����Ŷ�ݪ�>��6�xK���)h]jQ����E@�qY�a�m]t^�qp�f��Q�-��o����M|��#����{��9S/I�C���i���.��D�9�bͲ�h��q���J���{=�?���=��K3}��~]vv�WM1�'���N�9�K�?�������g뫺��jF\m.;�壩�N,2>YI4t�6�l�z�b0�gޙjs�A���4����#��^I=�p'��ӂFL���{_.�xϦZ�PB�b/�&������Т���8pt(f(���/�z�����#�*�ģ}C�8c:��,
oW)m�I6϶�~)/����
�n��+1��5T�������Rܬ�W��|�y)m�O	��M�0�ؠ�����R���N�a=�d��\��a|r�!U�r��=+04T���D��l��W�G�Q�}�K��G[g���C]����п��Fi�	j5�
��w���C��qOX��P�@��b&'w��1Ǆ�ﾧ2�/���d	/��S���-cY�����`�r�pu��x�����ۡ"�<ad���vT��BJ�n 2����|J�f�%lד��9[��~Т�<�� ���������0�Q��yQ/�yֳʭj![��q���p�YUNZ�0	��z.��A�u��g9������u���S�?��G�WS¦6(sw�����Q��^�qP�|�h�S�����Җ��6�D��{�>�SO�I�Y-p��&��ml3KE�{,��q�IW�]�U��({1��_~�Rc*�fpF�'ת�t�����'������7a�Ʈ�#�	��aI�;2���oi����o�w���yX�8�X m_2L$�?֜��w��2�C�ђSN-B|�މ-M_�f8�X��W��(�Y��xhԿAoe�+&t�����'-M��}!����c�a��Ph������6rJy����p��n�^'����kM�8딈��_JL���2�MV�a��������a#R�L~����W}ԉ��Gģն�����isV;l���4�A	�%��1�������4��Z����C;��tw�Y�
3�h��QS�VH��q��r[/�������0���Ʒ���9dg����W�r&�������%
��(�Rɵ����š�7�c�^ۺ�����8鴞�@dz,6�X��	�=�R/�Y;������v%v�/ԃ�����s3o�����<�*��%�͇��F��?����-v0 � ���.`����N�i��ס�~�ם�F�SDZS3��H�{�k`�»�aP�����'�{K���E�i���t�o��Bm���ߡ=�GD�ƱR�ͲֳA�eJ�:k�!aPHm�)\�#��4�0��������!z[��,Nj���^�! ���X��(^Gx~I� J��R�Re��1��K����_O�� �<u��@�c2�P�[q?�R���Q�ͥ d�ƭMİV��%9Ű�! ���m�Z)�s��Όa?=nX�m���xv�N��c8GfHz�a�=0 ѺYl��a@5F�����:ŷe���&����7Q��[�X'�w�n�&��%��M��_=���ןZ�j��;�ܸ��g6q��<t��^)����]��3_�{�V��8��3*`Ŋ��Cl#2�)x��h��m�~�ܺ��ې��6�M��m"Y)Fs�~�ن[+Yq~����&��8�]<�ޚsf�����1�J���Q��\�	]��&A/���Y��K��ō�Į�I�&��_��z��S�A��	�)��8�M��A��D&�0�)�t�m�e�s�%C$�VNTs�$YUXf�m�����P��J�)�'�cB��i��X��H�}��M��4��z�����x�)�$���j-W��Q�]Q(� �)�(6����s�0�ڞ���,A����a�š�7�D�\sH��nS��zw*���@N|� uM�84� ���K�♠�l��hfP�D�D��F���vʪ�U�#��"�,�"��}@��$tqh�KW8OEcźtч��ڐ���>,���A��U5{����ᗸ$m��H��]�@ U�l�$ E`?_6������4��{�Z
�����]��V�(��}9��h��t^TÓ�o��B����=��*���*�n2Oc���V��|,�P��QχK���3��Ѫ�וd��Kr�[_XA��"�K�9���X�hAH���0���F�f�w�O���(Q%���rv^��wE���EY&��Z��}��3Qb�:N�D.�-%B2���F�@q�Rֲ�'��j�$��y4sl�}V�_���E�lK��ޠ�Vӧ~�X��35ո�h�kؔ�l�j޿屉�v��C��\�m�"s��ܦzm�'���
9�ц
��,��A�v�7f�_b0��j�b`����9�d�Z�lC��	*v6�qA��ХF��j�}~a&���7՘�>���v˅�H/�
P�?9o�+�Ƕ�/��/7������� !L_�� �j&ぁo��[�҄f)�|�dPeL�0�7���oLǔa���	��@Z$���r�Y��~\����\"�z�8��3�\>+�<�H,�joi�Smv�B^�.��3�E��bΡ#�y��U肉Tϻ�UC���ٮ�[�U���� rpHٕ���t�v_�z�^�T���LDj�O$�<$	���S�:: d�Rܸ��zd��[|����1n�M+�A��S8��c���C3p����,Չ���7V�8�ә˰�h?�a��h�"|��C�~,|�zG-
�VR�5��{��k�����E,��ezzŲ	����rڬ�}2�sl�;�g*ܢ��|t�&@2A {zH�y��mg��
2�7*r��0~2X��m��z�o�JCi��M�i1�6�����99����
�?��C�� �I��M���YHP5�Ðz��#|mdK��'b$�|8#�Z���!��UA�W&"hc�(*��{T=�
�Gi�3�5XI�R���.Tf�{����9��*܉AF�������,�JXW=z�g�B�u�#q���Ta)�"��,�%�Y_#7�2L9*�3w/���}�WxX֞$�y$��π���|\�U6AR+��N����a��Eʫ+ wr$�������3!y,����M����?����<�5�qBɚ����P%t�VB�bq���Z�Ы�^���3�U�8�����v���ڿ�����[iX���Rձ���Ɨ<���P #eK7���.�������ǌ�j�Az'���0��Nhk�-�#e/bhW#�)UG�9���	���d�[|W�,���1f�7��q�Y�&�������U`��%v���_�2�����\��a����&�����pX�?OE�@�M��z,�wb�����0s�.9�T8��!Q}��5�Y��bﳵ&�և�Fi���aҠ���}��;�n�w
dʱE���!'a�b$�! �V��p�` �x�rCh���m�#��-X�[�Ӱ���*�I��>��� j����#1��n����-�i{Mz�ʌَ���j��z����i�>uSct�����ݩ�O0qֈቇ�C�qMI�(��v��ܷ-e���ʘ�ϐX	���~�XI���~Xjݺ8�A
�Urm�Ǹ�?��,�E&�	s��\��FfK2�is����;;g�L��v�Ny[RI
�?�����O�N�m��U_��dLVc	$[.���]v"��I���.5���;���/������o�7�C�`8��W� ��]|�*k]mn���*�S�q��\���K{���M'g��0�$�㿤�w�$� ]�n�W�sr��4�
��Iy2 F�G.6�ZY�����=�2�Io?g���T4t����޸�ߖ�m:� Hȅ8X�5�HQ �ґ1&fN�E��"���r���U���A�?u�h)�$���nii�SۨlI�N�f�@���Y ^W�Y�櫿��&�n�ߞ�^��$��0׮m�
�3'd��e���lk��⅁�M�l�C��`-?���2��6�G�W��0k���+�\��� ���B�/�g�?z>�I�f�@!}�E/�tsN�˄�/���v��-�x4��m�6���8�����V�_hd�X��&���|W!�R�X���T���'�m��.�A��q����P�)�T7-��_5:�H�������'��*./	|�L�N�_�"&@����N�A���3v�I+���.�J�W�aM��V%��=ν�cM�)�n�Ҥ���)+@D���k:�a�2{����ebh��oO�(TL�'���C�i�$	7�GcX��
� #Rr�ܐ4N���y����@��ٽ4�$J�3���LbH�����`@�a`	??J�ov��Cu�C�k�׈���/�w�M1�/C	2�{� $�0�7�Z���R:�|"��Ӓ�юz���
\Y~Ņ��/?����2�ر	I���ꄝ`��<��/v�e���*���2�
�ȶKU��E�P
��ijn�ҝ�3�g2�O~h�.9[I^�P<�d��E�?�����b�K9:#��	Tl!��C�K5��Gs@u���_���I�-6'u���l���![W�l,W��S�,��{._�����^��re�Z�5F��M�ρ##������X��5��IW.�_�\���-���]��N(	ǽ�t$B�DOr
.=��Yp�Ϥ�Tc}�/plY��������ϛ.G�غ�W�O\���VZ}�t+�p/�0�Sإn'arlMIfv�8�V�?L�%Zr`�-?��F�T4cc31��6����Ӗp�7���wrl��(D������}����z9��#&��nׂ�T$�^S3� �afU��i��H1-�flPBj�u�i ��~3��'����	p�a��G����Nּ��A�?	���OH�"��$B�;�Jv	�C�O�!\{QH���u�v�͉���,�0\�t9s$=⺞ji%��9l�� �ޕ��t'c�1��sP
��I�~=�J!,E�wm�J`��DG[ lg�}I���Ur��D=���SS��b�$����㚶�O��r�/a�x������
M�y�����x?}��i�/�o�D�^n7,�eE�i<�"���m�Z��y��=��R�d����׋�BU�<R�M�����>�CV�N��F@��#�4��vz���7*�f�m8�ps)l���/��!YZR+h�B�Ɂm��vg'@b�����
˺I�Zb:uS�t����i^*����;����O��&`�HZXꦻIO�e5��K�f�i]T4�\���@ !4R�"�e��E�|,#Lߤ)>���P/)��{\Rr�I��R`?{�D~w�����;y�Ӻǲ����d�!J+�3H�` ��3�WϪV�O�;�d);ն���F���'�N���q�uvz���vk���,�E��s��Hj�@mh��V@��`�vT��)����y�t>�1��ڏ?���:E\��@p�h<�?G�k���Vj����Љ�P�Yn�kKE�Avk⎪�u�����n�1;�72B�X��	�m�a�+D����	ҿ����e�?jw��|7���Ѷ�t�`�;9N�M�T�]~>�0��*�15<��nC�C����^Qj����3��F�����B2;h˘������v�Rg��|1^B�߱W��#�#��P�P����0;}Q��$"�..F� �b���eQ[���\���T�m�ѳ ��i�&�
��.Um�V:��n,�N�y}Yw4�&w�+nfA�?HbSӛv�
�o��/���z��r���ۧ���� �������7>UnV��k[h.Q��-�T���«��%mA�\��^������ S��W��%�k���4��&��p��\�[bt{	�$�Ib]8Jn�ag混y�d��y%�W2앚�_���K��"���F�)�ͯ6+����t���u�t�2.�&_�bnZ�ӋO�ϗ�%���1:���o,�}��Z������������C��d���	���pEty���D����s��\0��\�Ye/>�LD��_�����Iт�)�d�=�������4�}���v�1�+����Ju(�\g�n�L��+�m�ఘ�T�e�a,aG����L9��:��p�oX�=��*�w����5'�!ó�ԟ�$�#{S�Ms`e��[�_�T�X�H�� �"`��?eu�R-RWT@Z2����d%��8��|��W��D8 W��F�M�p�o@�B#/B��T��Ծs|;�q0S��cQ��rq.������	�.I��P���7TJ3�|�EJ�g�ǝH�+�h�o3.ӷ8_�x��~
!H���6�X��Å���tρ�MF(e.$>���^��z �&�Ï��|<�^KR�Y�M�oQ+��X�?(���ޖň~ڦ�bg�H$�,�o�%�[9�{U��x����vE�Vᴼ;#"����ˋ���h����Vyg��G�}dY�K�+5���w�Q�Qy
�<�|F��H��������T$�L�e6ʴ�t�$��t���2l#���:@�|j�H�����D���Vu��yI�s�+I��Y����Tsx��V�ϲ�	w�I\dX_i��Vk��̯U&�B�������#�8��f�)A�°��Ӽo�ռ^~��bg��I���Y��:�xƜ}����Y�4��D��ewuW`œ�Q��۹\��bH�K;w����p]��?H!@&z�"yM,��mg�m��̡�<o��|���4mE���$��$�a��|�ʤB�<̓2��2ro�W��Tm�%RH� x�l�}��~�u�_�H�0Y��a�Jv5��Jr���	V�!�È���
&��]ԛ�;�-"� �	u(��N �V���y���?.��*���j����E�HNW1��3nLt��)�wo\���t�-��L:s��q�J��Wg��o�[^�?Dô�z՗�2�.�t��@���1c~�DL��h˻����dۅ��r�:�w3&6��F2m���l&̓�(M�f�s�+C42���PSL�x'bI�U���c�u��O������P�+[0��g&�S�%u.��fyp�|>�<�xbQ'�4j0�.'�*r"i�_�D]
������[�S��I)��ך:a��j�Y����`�4:�b��j�^#�"��Q��uju�j�.| Wd0�;'DZ��A�xІ=k��`?� س
\'vH�)�qo`��W�G��/TvU�;�t��S��J����������D��gp̽�	;dP�M�a��*�*�Caռ^X'=�@�$l���P�z6���������t���)�f�`h_�����n�3��C��o�̹z�D���u���������m��ն��`{��̰��zN�h;�>�TG��T����fp��F���Z<1������A������9�`�:O�H_�#�t`=炓E��Nշ����;X�>�� <bT�K�����F�Oð�C	%AN/��h��"���Kn9�=����R��Q?�۞6�Sz��A�/�A�)��������/���;�ZN�w8m�r�B	d-7�(q��ۛP���^����k��P�V��J�]�{�y]�����*�ُ�S���S�����|�:K�%�=�����Pb�A�D @u�h��p���9��p��S�Ȩ�_ZAOv%�t��:����4�/r�'�Lb Kj\a���ʀ���{�ڟ��M�����	�w���Q�W9i��;���׳}�K�d%�:m�m������qv-�:d��B��a�r���=�i��=��x�a��^�J��y���n�����I��NK횺�*I(|��� �L<����S_����b���?���p�~,�]-�ˈE����Py��3�Ja���h��R�%F6Cm\F+�6�X��v��J9Ex�����#�PrD���>�hH�r�$9[=O����e!��W%�ƥJ~�T���	ɜ��N�jܲ1ف�Ce>+���	��q+ɘ.p����1�}4��P$D�G�e�i��Y5��3�����LjA��e�h���VM��2!"Т��G��p�!=[ןR>��tS�Ǯ��v�UG�ܶL�
��Lw�� �'A�J�s�c.N���m�'��`ݍN/?�{}�i�ó6,6�pɚ0�eXᙑj�$���TA���¹w�Lӳ��m���(���\7�3�?����C�|o��r��p����QD�(��4	�t� ���;�-|Q�P�\@���8�e�C�?� z,��`"Fa��6~�""%=�ݦAwb=��B�kX#$H\�[W��B^|�O�5�5�$��B� �ܣ���07��Fps�0�BcW95�q&��������DUop���'���P+��jZ�@�@ϼ#OE.��{q�y�|Oّ_Qs�~RvV/c���'Y�����zq�0�J��j�相Br����Q�|���R�#�����tf�	[!Is#	���4���@R�*�h���G��mz���q�H�_�ub�F�jfv��*��gt�TjL5����{�7��S2�F��eԨ���*����B�/�Pp'%ƸiFa���A9@|\I|�cW��#�3� ���&��b�����N��j�:؎V0o��K�^=ӑ�=������[��h�W�N�]Ī���Z�~���?�i���s��a��L�w����P�W'�Y ;k�����ce˙���g�M,]�.s+6�nE�&�1�P�;��K�z_	�0�(�m��Ү��yA.�lժw��x4�S�.1�ؘʱ�ɑĞ0*�2�Ha�vZsYKA���7/�$��P#簎���{r*���U�����^�*h�KiW��ܶ�dI��eG�9�B���0����>�d �?_� D����|��4ä�]��˻��3<�������X��L�{����6���O}�ȗ��n��Fn["�� P\��,/�}������ -Ϛ��q����� :��ު�$�S����U����g'���:��**D��
��5u�A�gަ l�l�vՆ#�/v�R8�LN�k�^t�J�?Kz�����Ԉڇ�n%}�afb����Y�w��W�B�B-J/��c�4��9hb��l���q�j�:_�+��"o��?R'�K,ܫa�� Q#�!g�t�W�H�E%�l[xe\ha����!�g����%��̳[�^�`�8)v�\�b�7W����w�#��� ���Ƶf��]�L��<�ȎO�G�,����]�|	9�<� ��%���{nA.������4^uJN5Z5��(��i�o��JO���1l�!�Z�J�B�F1���)F[de���o�Yz[>/�W~:!ٺd
|�S�n2ND:���A,�+�u�l0�s2/�&b@��QV�5H�n$�>:3$ě����<]E�^=��� ,LvVz��ƹ�x8k���D}��+�h	�	l��l���(��,�%LDI���������(����L�q�Ok�+�a�q�����>o�0M�J�`?�F��
���-�!��	�m�0fId�)�?�߶�a5�*j�d��j�Iv�$?0��ŀ�鲄�0��|J�`�^�Z�X��*�B�\��rg�`� �#��E-_0fLO�s�:��!��<��ʷ�CS�>�bD̬�*j�#>ζ4��7���\����E�qq���7�_��&�J=CA�ۮ�I��{#<���Z�v���F��@u795vG�F��z�����{�8Q��@��P�,���Τ�zN.�����*tVk0�G*�5���Nfa���A�r���z�?#j�r���M�{���Z@'��c_�61��o)a�^^�:冷�vP|���a�����J��=�Ĕ���ƫ����K�Fݲts�ea�!_˘S�MJ�����D_}H���Ώ�����[Dyv�E�����ɲj5{�5�P�}J)����Rt�<�����;
X�u����2�� MmH{��zGH��5"��$µ�"�k�D�H�V �W�v%�7�����?,X�i��	ͳ����R�F�d��:���(���.����-��`�2��4[4��2x�kO������W�zՊ|����'Q	?��&��qc���z�(<���p�S���R�f^�xC��~�ڟ&p�^�'�ohT,j#��]`��͸�(ix���8wt�vK[j�E��}�Vk�����I�`��'NX��=�i7�cݽ�.G�f/v���������y��bf�O��s�}����S%�n��"��|��R� 鋡A�]6�ӝ���f��BA�i��C	�a����`�U������-���*��5_Q6G���*	vo�}溌�?����ĤV1,��2��i���8���=x�}��H���y?y��ݹ'Հ2��Nq�"A�t%?1m�4�
���W41�����/�\�R>/tG�����D7��j�I�ʖ]���R��N��;O�n����j(�˦#��D|��L�.������v�-~���"^;$�O!� �s��$��_����A*��� �eд�jb�_�t }]��#�-�3��Me�����َGR\pv����o��q��о�n!�V�іic�a���O�ǒ�čE�?Z�H��y��e@���xS�t��R�=��Z�1������3
	�$R}�C�w[�qu���j
���B~	j
�-a9[`���:���;�I:9�e�5�a�TЈ*+t��������S�1+Hz�ev&׊�1G]�TE� )�6���%v }Y!�V'���;[1���36:����wf��Ƈ�C�ZHG��Yf�}�R��	ҏ�W*�m����z~�?4l��^�������!&�K��@����̮t��#����9�[�L��:�2v�7��[	�Xs�|�6�^�3�
˘x�R��Q��hYg�ۇ����'�"���~H��ϐJw����B~��ﵚ�{aD�m]�>�|$vC���z��z,�/{O�7	�粥�^ne��M�{P	� `����%�}�$��X�3�WJv��y`H��䓺�����*Z:��͉���"�;���c�L�B(<RS:����{�!f�iU9�k�Bnq��x��2���(�Rx���d�X�g�r ��/W���P	"#pesW�ԑ�WC��>��B�0Ң��/Ώ���d8��?-��di���"�Zi��O�F^�ØOR!y�6��6�&�|�D��v�YP�J�:��E��j���>���#3�]�?Ad��L��t��	d��3��A%	��l�t�2�+0�M����R�^K�fw� Q�����#D�r�sɑF�V�mRޟ:q����;Q�g� �(Gi
\����
;�%(�4�Z��"*����XxZ�6C��8][�х�ָ|G�;/�ղ��r?�W�xЏ@�C*�����\UB0s��n�t�]�XZ!�kr�z�%�k�g�X�,��jI���%�G�?Qs5��]-*R�����r�*��KJ�2a�����T3�Q�Bg�wl��3:���A�΢�m ��=>�.��w��d�.h�c9�d$ײ��E���#���\� Ė��&�W��>�|^�iR@���Â����EnN��D%�%�2��#q�lV�ZŮW�a�SI{��2��ϼ�5��5�s��|ʰ�bv�h�O볃�R�}򨉶��aU����&S��'�yw{��ē2�"��w �.w��О@1n\Ȁ�JD�����L0vՔ#�6ߛ��t�ޏgWz ~��eB���4a �k�ȧ���ͭ ^�)��i�&���L��.3���1B��0�5R�w+�Ҵ�&]��;}��)΂���l	��?���z�ʙ�M���r:5��I��*��qse��.k�:�E��0^�e��B�c\:�����%�5?��,"��"���a��
��^;��ȵ����N҉�~']�	d�q�,��އ�r/$�:���Q�i�}s���c�r	�D���4�����p.�����rV�v��}�]�Р1ڂ/����$��h��8z}΄��5����DY_Eګ���"�OP��# ]e�0l��*�8��[z�iMť���bώ�t&�cI(�;�c�k�k���W>�'c�R���N�Q�/��DHyGM�ۍ�t���^�Q3G�]�vy>�`��Eo\��/�Z���g���j��������lՔ_�_;���W\�s���q����"v�����8U5��ֿ'�س�Y���j�q"�d���i�#\^T�7�C��i-H�kO��=���_�zH]����^Ԋ2�}z[r.t@����䟑[��Q�&��kW���r�aVʓ�غ�Z.�qB��|+E�`%�뽞��P�ö�]N�o��sꎵ	�K�݀�X}�1�r�q%�� �s��O	|�Kt�5�z�/���犱�k����'d�d����0�ly|;ϴ	BÏ��>��J%�Y)�U�Ź�k�4�-qB>�>�Bお?�ʨ�����Lx�S&�D�&�a�S�ЎLL�iz�ϊA�%��A��h9�b+�Xb%W���w���w�zh_�_�vv:ا�J�əGMUTU��C��.�(�2ǨH�(��*T�$Ui#Τx�������<��$��h�~��Ź�:W A)�E�Um�K���e���85�@�)1Yw��ܠ&�$�&��Ee��v`ElR�j�)��ه�K��a�N�r���ǭ���ˑ&�!6��0����ރ�����餠��l}����#1�o����p�6v����1�i5�S�����)�́�Az+s{��f�6����H�r3-n� q4..���B/��������S���vxc_S~�ԝ�C�C~S
E��&������ҷ����9.�?�"��$���8VϬ��7�*�^��cdi��P��R��']�O�����z6u��'�p���m �W;sx6��0�vz��jΓ�3��v��hߘ6[-�f+�����߽�#��x�q����n�Tg:H�v��#ZFm����*�������4�μ���\Y�1����ۧ�RA4+�5���)���s?��E�[�����x�0����_���m
Ŏf j�I�6�si~��Xmܚ
xA�H6W^��=���c7��n&7���v*X����fDPV�	#�5�t���NT^a��O�//ѕo;�'W�s���9�;���F՘�bE0:NX�y�����b�ă"�7O�)��������F���S�����Ar	8���jK[!D ��K	ޫ���Wqqմmd��d�y�C�;�od� G�.���\�L(���^(�xHr����\q!��t��-�$��Z��w�B�5|�*��]
m�SxyY.u6#d?w�6<�WV�9{G�Z����6�3�*y�
�O�s>X�^$�٦FM䀧�Khx��]�z�� �V&ϨVZqJ
�Y[�K����bP�!�2D`��a�#��WG�������IH��>P��T���4�l@��AS
B����Ԓ�)�'#���� �~�P�^A�uT���&o�jN�W���\�6X=�\�B��cK\�ʻ����b�6N�,���u�}� _���ĽD{��@�9mP���}�/�v��gl��%k\�K?�� ���&��/���{x��H��f�)�A����0��`d�\�J�5Mߕ$QE����:�ػ2�9����u��3:�ђș�&/�W��lt��ɽнM��1�[�{S�����}���yA[A䲼�U8
#���
-����^'�A��a`D��2C�����%���F٩��Jߋ�(�5uPj'4��Hc��k��P��U�M#Z����έ}c�ɸt��s�b�[.(�}˲�ar]��I 5�@u�1�i o�+csK\"��d�Xq,��[�+�YV��Г��<�_\!���e�	���x[Bo7D�¼ܞ?����y�y�e"�����xw��O�����.����6�G2"�8߃{������b0��� �}�Ȝ����5$H�̴�<7iO�Bj�a��0ȽC#h����r�8y�'z[��y���u<��9���)j�*s����~a¦�+l�H��#)��x�~�jH�7�/2э��d7Ѱ��4�xgs����7����P��ɶ�QL�m���r��@k�H˫�Ѯ���g�!!R��x�SO�/���}F�[li�;�pm�3Ia������8�ヸA3�0�-R_-�3[ݘ�y��)���g�q����L�����0�L	d��2������M5DthQ7)3��=7M�	��Qp ����zB[aW�I����N��[_9):��ٲ�,�ln"��_���?�H����[Cu7�W�1\�Ct����7����Fī����a��X�Rk��4c'���Ϋ�W#���X<�|�HPcs��ã�11��+���ئ��WL�F��&���-Qs�W�~�ʦ� Y9EO=�+lBZq�4Ӵ^����� �+�K((��Jk����9����/��cg��}��2�ZM�K�&���#������$J��~�8���.�5+pmrv�x���S\�4��x�����	��ɴ�J ��ջ�/��Đ3�����O%�X禯:do���L��a:���Lhω��*!��Ub��5��3tPز��p�W�B\lI�*���6/Ȳ�D3����{B�:��E����(ŢŀI�"��L?d���V��rciFy�
gP�`5%������k��z޹.�S5h�f<�ƾ�V�Zս*�j�����`Z ���6���R�)Y���*jN3񋇐ɧ���j���t<�Mv����"��N�R��%벑Z�b�ɉt`ƤڥT�����iD|z���� � ����I2�
��`��wPc:��0}�=�T�;;Ra4$Z�	�IQ�K��"���O��z��z6�n��j��vҟ����S�o�`{��`N�)����׃�>|�+��|�m\�8h�^��N��+��5�������3 �݂F������H;�� �V�5���K�
�\�p�|N1~nm)�R� ��T_:pq�t����=�y��)�-��xܳ�ϥ���ю��Z�eV�)�=�Y��Հ�[c�rSL���P}��40�l�1Z�V�.-]u̠��K�G����F�4��[��l�sJӼC�g!#H���|�٬h[�2$�cL(��Ss���秥n�����������Y5��PƷ�]��5N��&�N+��vɨ�C�'�YTԩ�Mu�c�b���k�������Dnr�C���l:������*��o�1[�M�`����v0I��'�kF���,���6�ϒuX�n2/r�ޝ��;�*�Ap�Bȁ�؃�ۂ����[f�鴅��������N�Q���Lў
��1�N��B3e���%~�ͱe��s���0��&���S��Z�=p�x�|� ��H/��������հ�u�7�vJ�/��p�Q�6����11�"YhU��>���\������&#�ɷ�����t�!NhI���({OS��FA
���N"��o�����TG%$�:s��&��m�����&p٠�<���t`3�a��ߧ�̕���CQ5N\��M�l=E�����x|)��g����n��j��$y�1��.*C�8I�����;lX�D��Z��j�����-�<fU?ȃ�'��#-!���ӯa�?��~��,��f쎜�l�2]Z^��GY-�׮��s����Z=j$x��ɒ%�ݟ�� �3:�o�[��2�����0�ʽY�H;q��t\Ox�-���6��ʛ��8w���0_磧�> y�ޘ)�yľ|�t;���6WYOVu�u����ue)�&	� ����mT���8��f6�-��U�<�eYڀ�ۄ�(3y�Z�#��)�$0 �t�G_�R&��W�x�6�!J'��&����;�驞�sr�e"tf �3l
��$b��0��WM��/-���\c����2�o�@�����I��e5�Z�?�̮dǺx���x�>j�p�d�#�+��TF�s�
e������2#ӹf�>��Ӎ�T��u��R�]�[��m���Y$�V(�>�$���,�J���Nq�A�{[�f͌����c	n����*�&mi����|�~�q�nl���<��U�9pz�<�q>�i���d�͠��9YᏖ�p�8T�3]Ht,�(�����=b�����{�Q�ߜ����Ax'*.�wQ�T�n�?��`W�ׄ�l���]��)Ԥ'�N�A_���{��}:-,�&��*��m���a'�:Q`$��O3n���o�67c�T�0��`;s�͎�M;ȓ��>�7:Su��slS1ֵ�A*dl�?�@����q�L��������C�:9�AP���:Z(ά��	~�[G��k��y����3k�ܭ(���h�8.�r�6p����P$�j��Ҿ	���řL�)�R�%O|d%�G��"Փ�,O��1�W}�A)�K��祢��	v���H��;�ƒIu{m #K9��
-5SA�w&����?̴�k��êdʶ�&|/J���H�<$'��:e���ݗ�,�!��]�D��:x��dX~J�����t®��YR��'���?�@�H)`uEc¨�n�����Co}�KC��aqV5��6��Ա�����E��śd�wr�J�AW�ua��M^�\-��[�:��ݚQA�FXJ	� ����ه��!DKd���������8���%��0h�H�	�'�:�!��	  �ӏ0I������c���X]gV����7XT��%蛜�(��Y�+���w�I�\����guP��Yz'˕?��Y� ��F6W �÷ԧ����=hK�bW�7��XH�{�]���:�)c� ��|���?dn3S�.-E�\�$IX! �]x�%��6�T�F�Ip�f��q6�M���;�7��("���Bk�R=�v2�0w�'94O�nf9A~ŪC��_��zt�nS����V�����aC������5��,�)(��"��]�aш7�P��=Q��,�X��{����<��X�$�k�xf}17�m|���'hRH�e�U"���rE�u@.�Yʪ�|%��E���k2�y��枎+C�@�1B�w ����� țD� ��J9_����f�p(����(�Ls�����3��;PCM�H�>䍩,�K�.�kR8=2?{����)2Ci�d(r�@L[��jF��.�V��y��QY����L��#���o�y	6�XT�&|ĥE.S�셡tp��WV��;�F�Zji��<�l��a\v/���[Ǿ2��<����AA�]��3�y����{�*�y~&�p?��i˧1�a���?��`���ֵ�;��<�A|FK r*Z���g��QC��1��Ȩ&U0Z�ǅwu�!��5-�w2����;��pHӵU';<rb'�4i�X�SCi�{x�뿀q8{����ZGs^���"�&�ّ�_�puR�d�QWAف���n�@�lߪ�q�L�Z)'����Lg�΋0P;탴�}ï��Z,�'�4A9�q�DV�M_4N�����`������I������C\ۑ �a�����G�;atC⩙ �4I.]s:�Mȗq�5���1����¬:��WG50)�{7�j�A/���)��%��R���<eA�W�щ��F<�'Ɓa�L��Ĝ�Г��V�_�6 ��$z�2*����g�g�M�3@��QG����eвq�]�zb�z����$��;U!��V��ՠ�k	*�O��u:�,����ȓ0�%O��:��(��	C�ffu����?��/�(�F�������ך���:N��/L���.c��KD�e�"��9�sC|�+�������"�W���~����(R-�R%��*�!Sݭ����R�Ǻ��E�G4��Һ*�9����d¢y�9*C%���g��ܤ��G黹��h&ؘ�H�\�I\�'�����Bu�(p�-��SL��(��rٴ�v��O��&��l{� I�Za��6-)\��h��WxE?��Ґ��V��^"�D�u}�j�哘f�|
"��h����������x�b]P��Ȅ�9��Aq�)JB_x�t���h��ĉ��o$㰚	=����S5�v��;�U!�|Y����v$wZ�":-k˛���[&�Z��{����'g�묋���S_ �QK+~�C6���lT[̗&I��E=I�gP��_\m�Z�W~�����u%��?��	���1�U7?ݴ�ɋ���'M�{@m��8F���_V�)�R�_F�W�gd%
ou��>��a09����B+\�U�bwW��%U
��.:ф6T�o7�v��~�:�
iu�o��!�OĜ���d��=����ם'8�P����|�'O���Oo��49�
�mJ�W�|͛|�JxP�N�>�����Ge��0�g����-�I���W��� -d��%\�`���b�P�޼���_z��o�~ۮ4o��k>�`7Gro�I�	��r9.e�r#�(2�t�%:��i"�5ڪ����`q|��������=#�|i�`�d�}����:�;��8O����9դ�fyŞxw�=#"�ґ;��/��3�{����@j���ٴJ���hDq��_��v 1�.2�r��[���/�?���W���g5��ba)�$��#L����>�Okf�����Um/p�&�\O�d֑݋s��%zF�BpF�5��D���d��w�5�媳��~щ 5���ǁ
6e�����jK]�v[���K$J\���� ��.�-
[�1Ry>�[����s�{��[-�n��k����MYg��-ʼX� ЦbaKA�����e��	����I�S������Z����ֽl�d��v���A��bћ��XGw1�J����NE��f���Л��:=rǮ,~��D,��k"��r���*H�]E�M7	�(4(@u
V�\Mv��&���W�=���ٖ��%���8t�x�@���JL2�(��|�$X�r��[E	� ������@q���>��ރԚ��ͮ���ܫ��Y�0��M)���T�~"�{j)�%�^��1}Ҁ�%��y;����dY��e�E� �8�b����)#\d�Mk�i|xY���'b(懧�!�����W��g��|�=������ey������)(@����}���&���N�%�I��G���<jC5�|�ЈL�����%�w1� �Ƥ�qp�h��J��c��t��HDFxJ����
�Q����A��-ZF쒳�q?��ۥ����wE�7v��+X	nK�Ei:�M��^��we���(B_��a��Y�CU<��h��|
�>�em��W�����β�NQ�ju�i�테�����u���A�����p!�F?���@P>�}1����|=+��K��}��0��o<G�C��t����UHh�����{_Bd=�� +G��@�G�u �����F�Y�/�]�fAE<ũ2�M�H�O���^�Q3&ʯ����wi�t�Y|�_R��:,j��l�h{ ��%�	u�Km�x\�d��e~S��2����:�ӷ���Fee�_��b�)C����b���\�Q��iіo��.$w�Ɍ����f�n�%��$֖vw��C�XK��:u��&]8��4�Y{��n9nH�C��ȎY�;�Q����ȓ����&��6��������	o#� S!Q�\L�D@t�EvP����Y���$�9��0�V��s�) ��y|��ȉ����G��C���>Wm ��YU���B��;L�E��`���"C81A�sk�a��U��2�AE��l�fv,hG܆L�V�����^��t<�}Z0��_F6�>�~������b�q�b��6�+�|�U�p�J��`���+��I��|�#N����W֌�_��m���7C���[|�����C�C;��f��~H\s	?c�S�L ���xX������j��LV)�������h���*pfR�q�\�$HմY�?�vPG�!,��o��� �%��7 I#P������eƴ���"���0�:;���)0�)i�}����`{e>f�!젧�z ��`
��`�O�!U�{��6]�c���ّ8M������M����.Lҙ �_�F�`>�a�����8�w�L\hU�%���{�﫾�O{|�H�
�=婩��23ȅ�&3^�>�O,f�!�r�6<^��Ō RCX[7?֟��6OŇ�>V�1��0�t� 曎K���(��ǳJ�Xw�5U�ҿg2.��Ȧ!�Su�Y��E,H%��(B�;�P(�� =�Ime	&�vr�H+Ek�==@�ghπ/�ņ�ڙ��^���E3wxeS��	��"�ߵC/�W�Yb���5�ht^��W{FΧ��:�b�M}�*��hJ&��6��^R��fMuV2�>i���O%�������������������3
�)�b��$}���Ja2y�����U��pxj	�hVx��3҂�����N���K �2� r�)x�#W&?/�~�~Wd�0+��b�^�YdA5�|,"�ʄ�CT�u���:ܵYΆT���E����,�	F��$>ܳ��~�^KIZ�	�gV�;Zbs��-���YVs��Zs̄5F���A��}bjۭ����ߚ�Mi�p�1z���H�#�����(G�N�)��z��;o�!ݭi�NOg���%���$(4~��ͅk>Sx&��H�qA�h"|m-����Pܴ�7����t��Ǚ��6R7S��mz��;+��ji0W[w�T�B *"���W=%m�^䴣���&�s��`--���}��ys�6<zH��<�����O��S%��OC]�����As�#��.a��V�u3�%r�EQ��m%�9oW��)ل��3K��r����caw7����{��7H���c�Y��Y���Л"�SY3Q����N<;@�*Fj@�!���d�a��z&'������q��<�ӄOu�����J%ٲS��;{�V�|��◕��*K$S2��*�܍��rc �������q}�UE��N`��#����>�y8rT��2P8S3�S_X��{v��*��W�ףuzݟ�M��6�L �/wW�i!��
�|Y����БKspQBB�e�#b��T�'����Y/k�C���w[w�����3�C���ϔ�P�3����lI���!B��[5�/d�y���9�G�J�,�-z*`8ֳ�|>�_���A���c+rz3������Y'9����n���Pj\�/jzq�w��w��/�\�E�a�l��N��qT�.��.�[����Kl��m���䙉�,OY
݌in��t�����PIJȘ��,{�����D�)��Z�1�aL�oW����r���Y�ԫ�o�R9��
��������/{��&	�b��"L ���P��)�l�|������N�z���ǃn	_dO�B�]��;���O��'�J��hA{��N�����E�����87^2�3�3Eݗ�����֊�0� @�DF`�%�ĭ�x-��V�/+�/�HS7�EbgW�kNN �����`˔D�'�jk�L-q�V���9]4���}�d��D��-}�^pt�!(��9��[��ӮU
/��%�B��F�ݘ��ԟ��C���gQ�aJ������s6�I3с)�����,�p]��x�%RK��}�4��W9KzE-j�h�w�	��Z�+�i�{��§�gx�58`��4�x��M�~���~�(քj�YO��M�Bz}>~0��<~ę�s���:��~1�K����8泀�]�D-UˑZ��'R�a� B�0�}0�r.l;Dm����.�9H�>���	�	yl��Tz"�/��.@����l�;�d���8�n�?�����nHAWs_[��3�m&�"D"���5���V���z��.��N;������>g?O�e��y�*Z�tV��%߸��I�;`2�9���J'O[^`�S�fn;��`)����ͣJY
ړ㉪$`Y�Em�5)���k�SS4�9Y�����cd���+w��s�	�
���q&4�����T5����/��'�2���I��PI��!�\Hki�~�)?^���A��?؁^?���?s}6K����?�J��v�K�Xb��R��ݻl����ǄD�|��8l�yndy����f�|�>{1����YzM�.ǆ��(w�N�X���>�I�rJ�6Ml��$O���r\Q�@�DL(��V�T�[�!�^j�B���4��N��֚�X�ٱ��y0�֦
�}zlެ�0m�ޭS[b^GE��h�J1�H�_ ��ک��ffx5�
>�u�,��-�˅���_��/KJ��|g�W|���ك�����s;����h�k���m2�8)�_ʮ&�@x��� =���3���(�{>��՗ه���^.���+9`����S|���B��O4=�:�-�"Z��j*e�#a�nP3���M����z��>l�����+.H�4�#����p��D  7�!B�\�}>+>Ձ��g4!{(��|=�5��"3)�~�$_�7���Y���O�%��	x�_ ���X��=��LŢ����Z&9�{G�F��do�x9���;Zְx�=>͑?�>��CW���O���'��/�	����> ���/�:zȸ��a�ϱo0��N�H�E86���s�pu�1t=r~��F؀�AI��䜌΁[ �t�*,����BF�<i@����Z.9D��o��q���%�=�HOM���O�o��Ρj5\�&SA��fz����I�<Y�D�=A��"S@��b�YK+���uh]�("�:����߈
�٬$��L�
lT�=���읂�IMB]"�t�R� ���O�V�T;s�ㆦ(V�霄xEO!O���n3�̉�_m��v+Q�I0��O޷��M4	��X��Rk���|�\�R�_)��_8�KU[�5�#�[�o5B�:�������+��s��O�6��VL0*�0/}d?>�V���ɶX{��Zo��X�׽�)�xH�Qg5��ݪ�#���ߝ
����;�4
�� ���b��#@1>��0D{�_� �/�;��Y��Z��r�}��NN{9~����6�rT3ޣ#s�R��U*Bh�p3�S��@"���IuE|V��)��U��������@���q���Ì��é.��B�<�=���9��u?�a%<C"iցk S���0�⬒��	�t6�B�]c�-�VV�æϡ���;�lo�7�!�h֋4_�}�����P�@ܫ3ĵ��X�7��D�d�L�i�4�����ό�l��40�MҞ�$Ns��>�d�J��`����c�u6i�h81��C8�%E|��8«K6�`m�V
���
�̔�jy;�1]	����X��@��-X�����Hn���3��G���)�w�H����2����{���s��ݎ��*����]��)�|-�i�͍�U���7 T
��U~9�� J���G #�ͪ&��U��jQ�V ��U��4	�+;���~����O���m�y�32��O���2p�wx��#�}�2՜�U�]v��Z���5����G@�:����ޒ�uW���X�c���$�J�w��%^�r
2V�4m�6���Y����J�0m���j�\z��C���}�R�L�=X���_�B�ӻ�Jt�b��70��1G���;8,�l��{X5xL�@��<ڤ:q?�OY!����ժ����_��/T�ge!4�_������o��^�)�R���'i�u�8cO�c�$U��Sq�]�EI"�a�L\g��@�Z6�zJ��r�����f$xw��J

1�KM��"r����A��{m�k�?���ꆲټEmRn@�mJ�rA7'�O>DX{Ƙ�Ҍ���ց$�tg��n�P�|��(RflN=)����&�S6��f��>B� �t��	�f���F��K�i?��$/���p�?G:���<_��<A&��>7�b�3)Ga���'��8,�Y�|��֪�Ů�'%�������@�ׂ&��V������_J�'F���� 6�i��t�ǅ����g�ј���W��%!�^%��2 ��%w�gEǝ�H�ݨSv�`C�*\�� �J �>�Ƽ���h�q/V����%���zυ�Q�#P�r^l�]���&������y�0���r1I6�#ľf�h����-��vV��E���Uw�g���<Ж�^��d�iݹ���)Ý��T�F�\x�$(t�ǡ۬8V�?T4�&��ʌl��yv�@�e�T��{=:�������>�V�C� Ď��Ε�	rpl0��#[m��W�bU�~A�����ȥ��y�~��1|�ڐ�M��9���VDhP������&tDŹ���oTt���[U��1�AG� �V}Ox@p�29�2>�M�-Ƥ�a��	˧$��g5M;)��{]"t�P��?(�yf��(J�{���1ͺ[HT7D�5��[�G�Ji�^?��H�	�n�_~j�s�BL�LX�C2��aR8�̛�`լ� xW�S烇aC��k��|�^!w�k�{��Xb��o��MV� �`���r���v)���O��Iⷴi0-�o�^h���!�#x��]*y#��8�j���&\8{�1����<��:�z��|��.�l�R��R�9xD��.�˴ C�y�͆�}!:S�6�{�E�x(6�ų�Y���y�#�itP��d�4�۝+]���G���&0Ƒ�'?m��������,>��������E��F&"2������)�^8ԍ��^�B�H�9�Ȁ��f(��v�D�(�"��&}����������&���s�Uc0�#{��'z0��iϚ�(4�T'9|h%��U�W#�U�{�D���8W(0��V62�`�vB�~&�Đ�R_�!�Ȅl��8�O�D��_V� �[�P�x���ʶ�"U���磝&Fl�x6�l�e&�0* q"�	4�FR�[���9�ͮ�Da�F~YuK��I��bRB�s�W�k3-��1���%@2u���~'�"�D+9���#gDaj��7������1������(ǒ�p���۩���n����x e]���~.%uZu�pp����Լ���<'T�ߖui|�_'2ᢾ��JP���-!��ɛ:UHRҼ8�ܜ��#�vt��j��;��{��/�9R�*���ɋ��Y��S��՚93�ފ<�J���N2Sp���@�#����=f2�5ƯR-60�&/ST:�jK{/����[����ޮ��Z�C���8)��3;ᮙR�]�/gkJ?a��Y�&h���Lo�y����].}��K���Kd ��08�g���bk*�>�g��B�tAbw�JP0t5��̨��i�/�3��i�#��*�f}je~z��L����>$��٤e�P�/4E�"�ހ��`:s�z�	+���b�)<��"I��Y�a��P�^�Xa���^ Ł��%w(X{��~�!��L�j5)�0.2�_�o���eq&R;��#�_�X��������[�@S�j�.���2��nqC�7�7���Y�IѪa�q���ئE�_���-��!O���Bm��q*t嬣�G{^�D�c��ڂ�|��3����9��$�W(�kT�X��Hj����^��{��Q%u-Yk}�A?����*�n$[�JEE�ZJq&B��PO�2F�x(�_Y
��i-t�f#\��`m�dr�,h��X��<wb��-��ԓV���(^v�b
}�=L�:���R�T�
�Kd���%�� Y�	k�(��"S�luìb��;��o��&���Y!oj��?�\b!�P���5o��D<��ʂ�������j�?�?~h�&m�0t�*�fy���mſ��K(�9�����C�	jO�a*i9���u��s`pK^O���Z_�v�\�$A��V�%��l&��x`��#8��"м�Xx� �!�缤ý�a5���E�ܘ7R�3�f��)A�L/ᩥ��	@4�"�ܣr�����õ �l��W򛐛��.���C��Ι�s�WE郹���{h����k�ˮ\�ID��K��.,`�*F��[��
�� ��/M�J�����t~\?����	DߏN�=[.K�	�(�Y�[�Y����0�|�����r?���2yP�L�]<���ܥ�kɦ/B9�7�|5�鱎Zp'�����/1#A�[]�s�ċn��'�|���3�����5�nؾ��T����/h,��,�|�����&Y2��/!�J�"�a|ͮ5�ǞGw�ѣ�B�D�m$mm����!���!�Ktw�q����]�(X�W�L�����H�����a���x��x�@@ϔ�u3E5�����������F�B�=� �V�1Tz�a����o�Ir>ƎpkEY��Nuo�\i��3����J���OL���h����k,��~�z�kE�6�H��(�G��$7�����W����������dWQg�*�bz��h��#�<�e�l��d���A"Ӕbf��@���6+���{ju���P1}P@�¬r�g"��T�{�����:�T�WeV������`c�M'����J����;�]A|�>�h2�L�u���~�,vN0��������(L����a�F��l�Q� ��~�Gy-�[
���w9�#{3���*1���e�[ų����|I�Ɛ��B��u���Y�SHᘏg<���o�遟m�e	a�mufN�^o�@�����X-�D�m#�ᮼw~mנs�Ӝ�/x����
g2�s2�d�Y�{���zYt��PB���9`�U�:G5&�`�iCvk8��r�X�*�%��}8��7�[�,�7��,�p%>IA͒�T�����2�2Ch���Rض��ez�:�ϵ��q�(A�����Z�`T,o��m-C;�t�D�f�#���������Ux-��m���e�Rk�v�o$Ss=�ב6�Dяw!d��7������}ʲ�V	z4[7�.���}�f�,LEer��)8!��E����OJcd�q(3"f�"l��G	�;H,�eGѷZ��U�C�I:mK4�����9k�k���ίd�d���1��_m�=rʣd5UT�h�鲘�M�h��S�(}�)iѕ!�~v3��W���]7�2f�`�D�#�0(7H�J�]I2��7<s|���EZ����j<X<�2Q�HD_dB��j[ߥ���]/���~�(��ʧJb��Ca,��� k�Q�-Q�-��$��`�@�!�x���w����=�F�<|>U��q�Qb{8����a�H'���kV�T�`zv��6��䡈��H?��?'�5$� ͓�c�hࡠ2�]�v/�Si	�Wr�hA��~nIs�<�������Z�	 ?�o����Td��C�=L���o�t�[B��#"i�U
^��l	����P�@�"��J�Cm�OT:W�N�j��	W/� �,GS�Y�pcg�]x�N�W�̢��/�X�by����>	����9#mn=�a7d=z��W
�w�{#Gn�+薭ج��ٰJN!΄��}�6b
&�)�e�%ŌP�����T{�l`�9��/�L��K@�a�Q� ���͛FKQ�f醸�,�"6��ڣ��R�4��54^K�m�%	�@j�bY� +^Qҿ�?v0B.��E�_��}��V�s2�eE!�4P���L��nĔ�:^���Y�`*r��-�	@�;�:�Ҩ$�Q�צ%I���2��n�bo8z�{Wz�RT��%<�7��l��ʛd���?�j�g��� a:�W6��D�R�Q$�*ؔ�*FL;%�1�JHn#����]v��̯��v����
��;��7�Xt��ﻫ=+��BՕHpLw����u]�Z���m4@��X,8�'k�q3����"�hO����k�u.�_�zv�ߍ.��^BQ�e&�h����V��"�&f2Ք�R�LDI)a�2�[�S�����~U^� ���0:�)�f���5�EZ�]�=|E�ץ{�Z���v�p���JL�/��fc�"Z��a,��:O�b"��kz�̈4=�q��o<b;��Y��jGWA>��Ml�&�U��揌���n �q�]��-'C��9��m���п_�>��Ƽ���+��s�Gi����A,�>}qC@Tq����\�zW����܈򉍵���V��a\�X]]�:-"l6�=C<l�'��~�B����3��s��}�b��C�tQ�w��KX�C�m֧������:��(=H^&j<8�9��nr&?�)>�q���7�}DH� -��F�G�2*����V�����l��E���Yc�q&���b����۞�Q���:*�mZM@�Q<~w�!��\w��E����|�ύ�ǘ�I��y��j�s�
~�r����g|�_ǎj1��z�����x=��q�A�cy�`��{"p�լt�.�Q�c�l��`�.HoKUڿ�[jL�J���ԓ>e>ɳ+7�]|3�J�� k���/�3_;e��t����O���m5Z-v)���tV�&Pe-��N(U�D y�r		gL�N|�hD�p�Ӏ�ҍM�3�=n>L$��������[
P5�j�a�-yI�����x��<�Xp15Ùi�����D�)��R����tqq���Ǳ�y k�_�2-Qy-P��#;��m��G�KDEjwM����m�U,b5��3�-;׶�s.�7�L�N;����"Z4׿��+�1eJ(֏�3��hk1�#|Ƀ�'��I@TC���#Y� KN��;�����Bu�T�x�<,���v&�_K��0$﫜��d�"r�M������+�FJ�Ϧ}0!a��ο1Ҧ'�o͜!6�h���E
_��T�V�K�&�h��N�a{�(�Q:�U���a��rYse/��Y�����\d�w#Ł���F�p`�����u"9����vX&���!�c)gh��?�g2��@±KPAH��ǰæl{6�.�I�j�o�������S����ܖ��׼_��Q�?%M5��	�x/�&Su4�&���5�
 �U��K�(#��y�$��o���T{}<xoSSI��.(��m��Y%��i�آ���[�,�q��xi.�R�.�����Iܺ���oc-�}�(1M B�G��a����;q9S*A:���/���N�����W-�r2s���*��))�Ol�D1�4����2��K¥��cR���Һ������;h͔�� ��jI��t�����lg$�y��!*��DBH7���������[�(s�;YW��f����@b�E��$�}�l7�9���0&�50��_�z����� ���Z+�$�ũq\�L�@�37R�}G���ֆ����('�̟�ͷ�5�򛾳:�@$ާ ��u����t�
�p��ErJ���ۢ{��C�\9�r�ݗ�q��� q������\	����&^�O;�~��'%]5���*n��-��&G����ƈ4r5�y�%9�=~�-�`��=A�'@��������I�L�㟸IP1Dd%��#��!.�Lf��1ri�5(����D��wXi4��b̕�W7���zBӋ��^0Ǽe�����h���l�� ��[v]�(|���-�Xݦo"�D�;:_~�>'��?M*�C�J�x.4�S���
�bI�]���?[�����r}�\A���Q]#̲�@��1!P� �l [���=�1�<MaԸ��>�C�"Gk�9��M�X���'k�t��;���4��Y�@A	�2�y��Q
\k�!߹�����B0��p�L�X�D�� ��U��_�Y��h��g!��i��:�D��LoSB���/���;��|i钐 3.O�*�<D�_^@9���4�{���R=Q�t����!r�g����b\��[m���i(w��u<��o�`}\�\��0.ˢ_����{7�~�>�4s<2�"tLb�+�[���V�.�t�2v4��'a����R��ՇJvfn~A�'��ŭ�@Q�{�~5�I�ę­g��2��>ܿ�]���W�\�RR�C{1��5�&�xgƯSJ��Mk�&{���?�K�mE�d��O_�\6_����Q9��_���]KK��S�80Dj3��7���dG�IC�%��#��Qh�e�N#m��X�JZ�.�0I�6����ahqau��N��/8���4�Tebk�������SXY��MI�	V�ca1�e��0�:�S؋X��B򧨯
�cVy�HK��B�!ЊΗ���~K@E���=�a�g�hJjY�����@�wC�y��'~=@�}K�-��yIĠ�+}Obb����K�K�"A�$ӗ���`Ue�Q�H��]�F��I� 0��r���_, \��2�Y�����F�Dh�d���3E�5�H��������(�ġ��'@v�`tb���`e��Ƒla��k@�uPt�|�`��j�Qfŧ[/+������k��l� ��p�n��xq��ɚ'm,��u�2f% �Z�����B�^]<Q[`�<S�G��Jl&�1g��G�DH5�_|*G�s�a�7��m(�NB~|�C��w��Iw��@AxQ�u=(Q|"@9 K���Jht!<VKY��W������m�6n1�ty�B�����ͼ{!�9�3kyۏP��b���hNg]��D�B/��)}�b�-;ITz�����ǝ�c�$�{�Y�0����5�8m����kNbv�շ:��6K��o'P4m�����_��W��=���AT�� 7��o:��a5��~0��9���㡣Ͷ�;_ k ދ�L��}YЧ#t��XZ���r�
ـD�E�@Y�o+�?�3֌"�!���,v)����+�A3\��n�F�}ͪ��+:�b��S�6
����;�{������r�ɇ�V^��oVk���M�X2��z�T8V;m�O l��JJ��}l������H����\b�TƼ[������YRd�����[W�i�y��0�ER^���$1G�|4������ �<`��L&�K"�^{���� P~)�Pr>|k�D���*��D�ub��l�96c�S���!z�h��}�#<>u�C"B�a���.f���$(�eb{pVɱZ>t}��wN~`n�����*��lC�oV���k�]K�'� s���i6���ߗ|�g�U��T��S�Ŝ��e3&�d�����4�;g2	��-P���.���sF3<z#%i�a�=d��i~�œf���z��|�����	'ѝ����=��d��(��8)���;uΐ�m�%�ڔ���P��_�����S����cQ/�+��!��H�o���5gX-��HVĮ�eqJ���>v~#�u�g��n�c���7�'�Σ�Om������y�/(���8;�*&����<I)̽ٿJ(��ީt9`._">�d�r��h���?@|HSrp�秨�z��fD<�t�`i��� 爎��]^a�4������Y�IT~�Ht�"�q�� N�ޫ���F�]��kCs���8�!.^�	����q�(�A,��,�Ӭs�����%}Y���g���8�&��4��j����X���c����M兩ݽ��QE�6[G�]_+E�b�?�+�m�ǯ��30�3xW>��$}�ӛA矇x�6 �4�.�q~�C�����i �!����`r�EHN&~7�[3v�1��ʯ�3U�x�rԑ��;tR]7xa��N��9�� ���SB<
�IP���ϰ3c��Y�B�8��ˮ��]F
l��|�r��f��v9Gd�Cl�ukf��qK�kd��	�P�ׄ�X���XBZ*7F�5�4���5�9�XWI�����\J����!/�A���.��ϓ�l�KD�f�(��v��0��=�l� ��4Xq��b}������d֛�|z&v����Ѻ�ѣ�V�J؊�P����X��S�}�b�&j�_{H��W_V���i�oű�δ#7M�vb(���/G_���=���������u�W���e��5�
�v��λb�p����������7���	 Տ'��8R�,�	_���M`������JD��*����r�V�۟��'�l�'�<|�<�F?1'8Dr1g3yX�	|G:X��a9/�OX��a�(˜"d!wU�ࠎˡ�$W4�7U2�mc=�^��-��3��uo�^Ԟ)��V�(͡`�s�Ѯ��i!R����K~UR�C�W"y������8:(��_7�{�d5P4NR�J�IMo�7p!U���Q�4>�!@�O���̀=]wT���je����5I A�r9}v�emN��x;c\�iG�8����@�L�"]
�v�V�vtiԝ��g����6���oJ�2��_!��?&�@T��T�����[;���9�kfQ&ׇ���� �
d��\:�x!�����P00`f{�X��(h	������dh��.��M,���iHי9A0	b�+���>e	���Ys��K9� ��N)�ɝ<D�F`C������Ep���1	��C�K4�'���h��̟�1�,�3��;/�u7ͣo�����f��P�9����Ґ�:@q�����S���cs��:�eC�L]��0�)}e� ʂ��O�Cs�d�	�e�x��$[���l��§ڦX���Ff�]�%u|*[h�i�j��9ۘV��߭<����<!!~Xs>�u4;��V�W��==I)G�:�D�{z����f><!Y'��b�pB�?��WEz����Go�M֕S����N`��+�^�fmԌ����-i�Nڥ���A��7�����)ہh�!��M�Z,�ͣ�� A�4'E���"F�5�1*'U���5@#��	�R�7�Eb�ݱJ=��%(
���
j�E^$<q��������h_S&�ִ
*����!^�/��y��Q�����O<`	��F	��e�p�T�2|V<<v��TY������������%WN�_Da ��yf	����-_�,<!<�/�\�J����PIo����G���9l4�ȿ��[�R=6_ϲ;@�UU�ulɸA��ysؾt}ıۤgp�q���K8#��|��Y8����c�!�l�xw: ��F�@.oy����b|U��j��7�����uِ��JU��n�K��kU��E���d�	�i��0�	�A �`�wKn��B�{��ݠ�L婅�D*x�����<���0��JFٻi�;�\�B�{;q�'~��X���/��ux����Fƥ?�{�Qy�#��R.v1�\�'�hf�rڮo)LUv$�fрL`��hL^;���P�{l���^io�E?̵��н����n�����G����������4n�Q������O�*Hq�����8c�"�ȇ��k����j4� ��98E"9I>#���׈����}̦�(/_TL䍠棘\�C�te�=�;˺����V\��7���Ai�+�1迺֍�x��_����4bo)�z��OP@�$u�����&kF��r�Ǐމ����>��!z�ͿJr��՛�ho16B�捰��Wz���C1�!p���P�FD�g�O)v��v��g
���:!����w�U"�)�a�m(J7�Q�E�9�� >n���/sq��T{mM�$÷�q,�͖+�A=�͡�;���������.�]��1hp�"�@��U��_�!|��z����m�I��b�b'x���zw�P|u�-�*�h��N��no��b�,��fޞ�'���_�>��*g-��?�T��Vq��R��*K���"~��]}Q�`X6VSL����0��=�H#36���-c���rw�8�M�BN��w���Z���t���`�[�����Msg��B���S��e_AhlI/�q���S��!7��ZA��k�p m|���"A��,���;��e��<�,�*T�Ġ,mR%;g)�]�|���qB�Z̒�(�gk��Gȡ��n'Gg�3��@��$1Q������oWv�D�ə��dK���	����#�vu^��+[�/��� �l�B�wm�v�@2cU�V�]l_f[��RK���͋n,Yq�5a�B�B�A��>�ooS�v��
t,���[�3�p����r$-ʴ�i(�R'D�^Y�4Gj�U�Θr�������$�T�&���z�l����*P]��G�r�0����jZ�@��	{�>5�N���Ā������nݔ5Kv~��`��Qj0�6J���J߯᫽%⟖~��i�3-�I �܉q��ZT&cM�mAL}Ź�酚c��|)r�5���h�c7�젴eی�{v������;�QĝՅ}��*ö��'�g���ώ��ҮC�x[hu�F�-�Z�[u6<X�Z���:}�z��┿�y�|�lc�e�(� u�hi��LA�zJ��_��P�B~�^A���Q�	��g:Dt��4�jƂ��E9;n@0c�~ɔ��!����a��cN��	��뻤B{����4��j���
UF��SH�2]���O�g7�\L����o� *>3fMl!l�kfq��r����;��Ě��cN\�o�:���:Z Ј�����DoO�|!Ձ�r����h������l\2�9�2�{���Ӎ,H!z7��ul�>����	I\�L��X�~��$.8y�7�[ã/��}�P��70�B��y�� ���y}�Jį~2��r�;3�k���*�Ҙ�?^SYp�{9�]4p�o�:~���	[�t��"�6f.29�"b���Ȃ`r(�s�0�Z�V���Y���ܴ9���؂#��9J�F&dɡ1F�/+�����@*aȓ:�3��#��8^��.�����W��fsȹw��}��y���<�O��`WI�d��9�䳤��3õI���s��L��і�����&?e�1ɰ�;$ý���͜,(=`�ݺE6V{��5Cs�W�zM�[�	����?�|d��9���g�U�O�E\�&�V�����m�i��M�R�X!��07��b'����xmq�/
v�AN-�Į�)\ҚH�nu�Q�������5�nꇺ����//���.+�.��&�+Z�e ���sZ�m?Ǆ��$���'�|�_.�8^a�[�N0�3��O��q� #���ǂ�}�pb3�*wv��,}5@�|E��#��$.�YB|��ͷ��<�,M������Z@<�)m�Ը�e6t�aLRv!"m�M�+|��YǶ�P��7�Y�O�uj��5*^E3w��K�̓�ZnGڱ|�D�J!�<����oh�I���1�y�U�:T,,�8�2��k�]._�9���4Z~�1Y��lԳ�+���@����J�P����I���#��+*��S��o�? Gs�Ug�������f�J�I	�K +�K$�Nl����&��2/`-�jޜ�h�<�1I�U�s8��)�;�^��@�>{�<i�ۼys.k�����m9~!ח�$p��[P�*���,����+Bt�(�l�,Ld�`$�G�;��ym�C��D�'v434��f���` D�)\t�����j��7�����}<� M)4�NS?T²~O�咕]zP����a��HʄG�JZ����_���Ͷ���&DQ��H�9�_�K'C�ߔZ���cr�����št.*����%Z@��٣�sKd0!���x�t�=�!��%Z���s=�����9�W^z�K�66B�P� �����)t�=�r����5GZc	�K���uV1|Q4��&�����
O]��g�K�9�<��r�s�g�G30���Vz�V糲��$����������E�|G&��HIS\vy�ِx�����!@�O��q���W��_�aT��y	��bJL���"sd;M`y�������'(.���9���粼���ص��{�+M�e�K��z��p�h��)>W���޸e$�����*ТT��r��}�# ��k�7O�MOX�A���/7$�X�����~���f+uΤ�!�g\�<������K���t�[�,@T�+JF�>��K��Sci[�g���Q;�݁�����>��R(d̩������ѽ9�3v�h�[�����Y�yf;��9���&��`^�6�7���Q ��2~A�����	=��#O�Vk3P��cX<��U��Zxg^y�aVL�Vow$��ѬN�w��C���^����3G������<���1��a:A���C����P��h.9�vr^��L��*r���v�7n��R��c�(l!�&B�ԙR�*����6+��;ł�IA]T��Kn8й��S�ӑ���נ|ݥB�ɵ�#�S�*�U�W>�H�W�ͣ�.�TK��~}�"�M<!M��x�՟�^�'����q�ֲ�4Lq���W僧�����i��z�8�ǊH�z�mmk<�UiS��%�v�Ѭ�v)J�+��C�Ñ�y(Z������(��#C�gZ���w	�:$��?i|F6�IR�����[y����˖_��-�2���zf*ں��3Y��Ng0�e7���Kbi�C��F
l�;��XBR�_�e��퇳$d�I ��i�F�4q��o��{l�#�<
Hм��)�?Y�˕�W��Wd�����CQ�\	���Ph���ac��B^�~�q����n;<��5��ֹV������Y�:�Т4�!���BlCyٿg��dK|K��^�(�Ib��ZX�f����o���61����Ơ���������$~�4��
�5K�ʞ�ߕ�8�|g�����T�,Wغ���`p�Y��\���V�h.3V �r�6^��3՞^�½���¸�ԨYyXk\��Dd�'�=}y/u=�N��;�d��A���7o��M7H�},�޶�4U8$�NΜ�F���O���&Db3�	�*�Dą��jS�iNs��cW���s2����Q.ϴcǉ� $IQeJc�vi\Ѵ� 2b㒱1G�w6e?�*[�-1�F}(�^I=F>��~7��;�8&�rb�����ZW�������ci`=I��Lp�q[���m�}UvBg�։���֡Ks�3:�5$�+�e2a���'�b��a$�*���\������[뫉���a��������sI�-e��m�f�e��a΢�U�K ��n����Z�Z��i^mk�ӆ��ѕ�K��|0s�aN'�Q%m��8��ntKN��_*�[1b��kٮ�)�Q�np�}��"'���7m�����t>@k���a���3K����Lo0�B�}��
���G��@Еx?�:ٹ��+������T]q`�V'j����f&�`��r�s��@D��d�v�ɯ����R�Ŭ*\o�;��c�MuL؝�m�	g�W���-E�?�y�y ����Y弉��Y��|�����d���u6C/X�nw�&����W� �|���SB�NņV��/B�Q���4�D�@���&�{�5��_s�[?�#���쿴b�/ iLN-HƔ�a�-m[7�SY��h�M$�q�N���FTgT����F% ��yp�{| ���p4`9E�<Q�<�p�K�#Ö-��Oj��pR��4;MA�p�����"9��ew��](�1�B�*�<Z�Kʊ�
s���'�Pr�J\X�Q�$���n_��?:w��݃g��1��,�w�mT[n>��	�@�[�*�o9�b�@��v\�-y�2ܝw:�e|ה�Ҹ��v�q�H$�}Zq"u�����Ge�5�=�-]$��vk�3Jk��.seu�6����I���^^!3+�(l�=߭��ؙ����ej9?�W��<��[��}�ش�1�at�&%,��otfwrM�4�lR��5(��5zg_vڕo�L���8���Z���,b���.8 ����	)~	�>a���n�U����}���aE�Y_�D���_���~灳W1uK��:�Ǯ��e� x9��&�8qڡ������"-ڊ��c;�3D�r# ;Jh;H�x��������$W�TGh�?*��5◉ٷ�DCb#���Vt������t{��w�k�W�f���h+h�B�#�G� �)���oܸ[�=ѡ��q5�
��R?�p<%}��Q� w�E`sz֡\�5�x&o�#@02�o?:{�x]V̅6�JkW�+̠{�RJl9��,��qָ>	E���2�;a�c���C�Z�_�Y�\�H����*�%�)���,˹)3�]CߙoPN<U@,�Bq�OM�s^�Z�j/���":��v����"y%�!��sQ˗�mf~��p�eL�c��A���yC�U�AO������Y��	[V�x�'D
��H����,����>wX9ێ��Ƀ��E�&�~�{�|�2�RpF�����\T�W�$�ٚ~�����e�yi�x���9����AH�2&3�B��U֚s����
i�ĳ�T�]�Nfc��f��Z��^��s��	uH,�����c�y�H�Ǽ0��x��#T���=R�H,�w��:	4F`4z���H����*d�����$cŠDQ:�"�.��⛋�R����U�k:�}_�;d��t�V�}����m�T�^���Į <��I��bF3O�ڔ,޿������mϯ��{����2W�UI^�%F&������CD���bЬm���.��B[�4�)�]���Td�_��� �7N�r��V�ʨ?�pm'�  ���,�����1��&R�K�����h~����a��:����s�S�A�u��|�)!!�$lOwC�X��k�n���ͶR� !�b#ު��Ⱦ�#�.����d�.�|P��Բ���\R��%��udR��0(#ǽ9PR[�*��"Yu��^�^�[����!��Z��e`���|��?
0��V��d[���ź6&�Wetk��$�@ƞ��¬'�}y"���єc�jɔxK��pm)А|g�W񇊳�	zuP�lywZ�\13F�-MЍ���ey�q���9K�P�Հ�N������x�n�׷#@����������?�i��Q��'��-,'�EL����g�WB�ս�����`4 Ă��E���v��M���}Vi�� ��a|�~���,v�we]��,����^��ҠN������sI��P
�ޯ~6��N�+fC��ߠ����LU�e�))���u�i'!�@��]W�@��ςt<oo��앰�����ʺ���%�B7Pr�>�2Z���v5�+}Fi��oҔ#��㩭	?���ٞ�Q�3�rX��M��S�m8���9~���xT�(�6{��ݏ,�(F��nV/���~��m%�ga��;C�<(q��:U_=n��W���Սdo\�Y�;�_��8Ц�s_N���)Aٜ@|<�w2��M&/�#��	���!>��6�i�uv�"���ҫ��H�^��a爇8�D+�-ڥ�k���T�g��H��S-�D�g��A�)��}'��$��ס�����?�8����-?���
Fk��-S[�Л4��,������x
^j�ڄ;����b=bٗ�v�rH&��#ase������ �'�s��+���t�l�HU{�b�P�`tU�E� $)��(]��%pU��w��f�a��T�6o����t6��V>��*�.�U���i��-�E�L�,�� 5~ujP�p���nVH85f���$�~���L[H����x���h���m���������# �h���M�t�Mіm�o+�P�f[��� ?ryV]d�������1Կ����ɹ4��u�Ȩ(�5W�$-A�R��쟋e�Ò����k*�;#5=��Q��l|J�h� �2a�%Oj�����6���d��GK��)y��PM�e�z�ā� �����6$�Z짒���@"�:u��Kj���_$V�h�z��?#Zj�	R�.���o�k3�i��U�X�d�Y.���_]�6����-sM�5�Z���W��'�16�j&��뿗�е�*PǍ�q�p�L,G�L�����*#0�Y�����tP�]�E2�0s�!Aa�C0k�c�W��yɸ�����ؒ��:F���c|7�˃��`[�A8���ɩ�(ߦ����QJ #�(�����z���|�/��t�}$kj9�� �w�>$��������O�rq �ٞzo�,�������~��-�)vJ�a8`^��8G��W����'��0Zt�g�q�(�x�V��q�^#���I��(��I��z}��|#��˗<�#�~82����~����L�ЀZэd�ۑRsY�L%�(S��s�>��$j��p���[��O/�m��y�B]�?r	�^%�p?�q���/�9��	vʻ�!E6fj�P3�ɭ�xlYL�8������^���O����F47�,���GX��cሚ�N�M��=`K��p�b��g=�~xD�	��|��Kz��v� Xj1E�a��L�(�i�2�6�r��@T(��2Mi�G��rl  x@Uk_U'�׆�� tC�,!��'weC\�_ֺ�&&��ƈ�����?���-Zh*���*l����q�hp��#�IbB6A�˿�X9�m�`�V0�Z�(��;�2%ָ�=^Z7����$.K���x�HAu<p�;�mϋﵓzzy��%�v���0Rj�=!�v��e�ȍ%me��G���w�mx �Z���C���L��NȈ�,��Uf�J!5�I^@�h(��ۅ�X��kK[@����B8iX=n���j.B�K't4:�
M��Zj�A`F2��9<�����+�k�0�eÂg;�C�\��Ȝފ���i�S��bh;=*@��j�|�a6���N�jw��u��;� ��8f�J�ڟ�n'Ġg���;y��]D�?qmd�`� �,v��r���$��y�@稍�V��}z)�8����$OJ��_�'x*-��]J�ݮ������B}�c���sM�J�*}��(���Ґl�븎t>rS��.7�`�������	ܳ�1�,��:��� D�<�h	� H�D [`lE+
��>��c�v�N��=�Zs���"i��ۈ*�>��_݄8H�U�8i�6�qd|,Z���0^!�O�;�7�}��������2o��f��.B'����A�����`����2�vg�%8=��m�iUu1�w��tP�*_�Y�@�	 Ĩq�2 w����U@#沞�9����!W6GJ���~�~���E,�JcNN��$���������R��}t�Sͫm|�7h#���fs��g�:��`�d+�&�����&�v��("�5;^���YgK��V{�Kb�W�[��rt�`߱�+{^�I�C�8j�K���%��ȍ�������C�[���Q�����+ٚM���PJ�'uI�fX�*��a4�"�)Gw�v�P- �!�;����3��"�.�mx�l(P#h�:#�)�����W� ���ʧ��5���v|_��o�W�""
|��̣K�COX���N�H�4�?�����ఽ`:�hD
'Q��Pj�8x�+im��$��`E�ER�>AQ�P�Ut���]������
��2ݼ��a��
1�K�9d�
l.(����p��+oo~z�j��҈8(�>nʖr\0�֣�G�2atW��^��1F|[��7'��n����D{��F���ٜ�����W�8�s!@���}Qv���e0��J��DY���-M��Nn��j~���d�>n8�/�B�p�t�l�XF�� Z�	+�c�'8� ا3%c�!�<�@
�?��4�(z+Rj_+��)JH4<��/�e,�k�75�U�Z��a���� ����B�k�4%OV~��:�H�n}�XXhf���FȊ�����O�m�Y�J�2P�;ļ��p��[
��H��vY1���lRc�@�7M���@@���3[S���4Ƀ��f�nwy��y#K����gB�>6�t=x��{��{�Q�s�ʃ���q��O�t�8d#� qgpȌ���(�O��d�1hy�fOv"�m��|4��N��ڨ�Ζ}I�2<��V�G����$�XV�"��r��nB��Q]��R�{�-q�T�u���T���N�ر�r����,����ܠ'��oBFV&e�z��v4�~���������uh�[�m �?ٗ�WYYpU{���?XY�.��椠�+3G�|cq����=X����g.B� �F�T��v"��X,�"�e���>���� �,:H�5�����BuuLu���EQ����'���M�#roU��ZE�)f���rg�*��޶��sSn��$��K��Ho�ELt�;�h��d�9�=iof�7H�>�y#̺|�֩���!�%Z�7c{��,ikN��פ���~i�"��/8�YJ��LЦ�֫.ݽ)���.�C8B\�X�Q*���m�<Ӯۢlߋ+է8�/��4���A1O��H���ڑ�!���l���'5Q�`629��,��Hޟ\f?�>y�sːx�aѨ�V3WD��o�ȶ�s�A��?D()�,��_�o�K�7���
��5b�]�l{�4OL�����2�̥.zI\��� �uc�S4S~ƨ�|�����<KP(� DlϺ�0�Yv������s]�C��G��+��u�$�G���z!�D�����n߭��(&_gw�������%����uYyV\�b-_�h7"'�#�	���s��-��) ����&[��3Xw�����z�+ʈ�k.mfB�T�*��r.Jh�Z��W��}&M[�䭪P��b�)j������N�c)���@+σ��DC7cZ�JlS�@��e@s69$n�y���]]iC�_�%�_�{��NL"��l�������s��Z�r+���ja�Qڻ�:�E��x����󝤫��J`ou=�3c�� �O���FJO�qT)�����.��D�����0��Pg����k���rD�1K�'�cG��rm�Z\jAp��^� ��*�\~�~,�a|r�eQ���*���P'�g��J�9x��d�~���0�թq��oF�`E;`��GkK��{lxXg�Y�=L���?�\�>��֒�]YS�r'��I���{�0��`�4�0�{�a���**G�}����E@,�d��U>�K�Anl�?ł�O7$F�H��-��e鲻uXc�����h��C����	y6��c�X��&R	GC��Wk�ohXH�p>����ƱT��Xx���ϰ�F�ȴ��}���DRw`�W^�����}H �0bD�b7�G?����x��|�a����?�.�F�����Y�vn�o�R�q�D�hE؈�u���:�!�R�)�wO~Qql[:��}���E��,L�}���uG��0ȭs׈��O
�Z
Iy���^��Đ�ͥ3֕�^B�{��W�w��Ԏ�pH��{�8��TZ!|bn�q�v�-+��b�VEۤ�S����+�ZJ�%{���2lg��%,d�6+��<������k���8��>Y��cGQ�V�A���B;"w ˎߺ ��1��C���ʒ;��H>1�._�H���]Am�!����s�������94��N���pP�w|��I\b������)�I�X 'd�͂�M��D����_�ɬ�� �`���zH���pn�z5���GhPb��c��rw�h�r")�+�pf�׼IѨ?��Gt��|ig��N� _����"�q�)U&����M��q�@;�e1�lX�*M:k�䝬0Q��术P�L��"ϧ�`���/�����K
M$xx��R���2�v}�l?3��A%rgJ"�����Lg���������n���dc-V��m<b��ޤEX��Z�F�3������n_�%�5�p���[�-��hzP��*	�ł�]!}�<�A�㟰
��P�c��X�m�C�����lA�� ��BP�g$�̙�O�ӕ�]Q}8-�d�d�z��+��:e���&����Ќ��OCM�*���5l8���Aa��`������v��;6�����?�#Pp�xK�^���H�sX0�.�����Xmڦ��`L�.�O;a���p��j�ṋ��L�$�У���d(E���ӔPlX3��9��իpV��8�'��Ƴi�k��;,pz�G���@�P�4�|�wFey������ؾ���J/L���tӷ<�::�Q4�H��~�۱É����4ۛU �E��Cb�i�6��������Ӈ䓹-j� swp.�kwv��E��W�y�����o�MO��?�>*Io�ӄ�Rd�"%�z�B���Oʋ�b�~�,~z�
}]��2�t��ܰhֈjXn�q'��B
�&�B��bX��ǉ�Rc��Qr.�!���"�p]P��Yf1���r�����f�Q�/�Hڳ��,F�Et[n��D���<��pSR>2$��%4��֐�R#M����T2h�l���z��26�����U�+dɡ= 9v�ԣ���u�#����ֶ'4��ө�,J+���!G��q��Ӆd��ؗ4h
|�}��l���8ȯ�����O�22ys�(��4��UD���| ?(�{���Y�!G�B����B�v��~L󆀱�gC�~����)V��+� ��ED�J�]�������u51{]'GČ�V��CS��w>��&���9F2j�A1%��Ӽ�M�G	m���C�� �I��ȭ�a���v��H7?!����H�IERr�"�U�Kx���Y����x)mؖ���J�.��|��V�(JJ[��}-:�o��AϜ�],�f�^�;���\ctq��x«�x�_�P2\�Z-C���t/��VR�� �M������7��sk�>�����t۝�m����;zK��険lK�]k~%�{�؁U������	F�.�������a��mhr�缉�w�N�_9�`��8� �7�(�s���)39F�-D�衍��:���#<�R�?�%���}֮޼�T2r;*<���BC�P�{�K�~�0�4���R��a�р������xБ������F��H%�v�``�D��7����pz�7Α�M�ڼ�h�{��.q\ѫ��<l=k��ŏ	�G&���î`E�],�>xw�����a��qT[�<���< �$��&�@��2Ny!t%���N�f:0W�����UY"١v'e�t���w.,���BL��.x��03�~��r�4��ǀ4���6�	��Q�s���]�H��vҫ����pA*N��1� [���Y`�xH2~�爎�$Xt���o�����9�W��Y����b���CF���g״�`�B��~��\���Q��ۈ߄��$E���9s}8txwBU$�-�6d�8�0�/�lT�$��o 7�j��`8lblce#c�VK^�SgTz��n�|@�B��U�dL�Y �.���q��"̗泃����6���e���/�ṹ��긾��a�GC�3����l9� o��V�lQ�`"��ث������@�)�O�s�w)8*8ׂm��ƿ �Xc����FL#���0�����-���߃�Ž�^�#�X��8������l3��O�(��ȅj̑C�?;���QL�pK�7�-ԩ�.���)���������B�:�����G�T�p�����(6#���3���M�@Ux��k�Z�2rFaS!�y�xn����cg�{)�m�GDp�\�T�`��B��ayTv"�ws���[Ȑm�"����T�j����^�J}��QD+׸��V��u�̩����Ϥa���k�Ƽݶ����j;��c�N���KYI0���ŷ��,���}lq������K��k���T=��@U���h�Ʒ┫�X��Ί<��6��ᶂ\�Yj_[�F񏜼z�7�~�-FѕI���2�Qù��5c-�ZxSL�/���[����)~	A�j��mcy�� ���U*tc�1�j��h:x��)c��DU"G·��7|��8r?)�R"M��o�l�қ�E�- ૙झ����}(]�� ê42ZOL�O�����SFq��wh `�ޤ�@�_qx c��D�m$��-����\t��g�����}���	�A�m!l�ku��H���ǟ'�n��âr����\�񄨞��Y�Q�v�Y�^��?z(<�y�X&0NȘMz��ZMD�F��p��b��)$'�aJ�7\��]	�m,֋Hb?0�/�+�	0g#����9wz��^G��䔂�P/�$�d�!�v"�>��<�-���3@��y(_"�!ݬ��Ozm޲��]3�>㤪���=!�`4$����(w҂[�V���[�^��"��}�[vέ+� @��g	���A�Z0�39�Ǥ��ꏀ�o�@�p/���I��W���\�k��x�bg%ѭ�@�R>�kr��(�{X�ی��M��sA>l[m�->H���Ak�L�J�Q �A�x�UZ�=��(8 9!X����y��Y(T�E���C׬P���ꔏ �/G#^��C�Q�
ȌD�JĒ��U��٥�;]�M�'�9�:q��%05���j�k9"x|�Q����@�^f���*k�qڻS�_�s˓T;�1��P�c|,(��V��B��(fzO�[6��!� Bjr��w� �Y�ي%�C� }c��	�p�;/��3�/8���j��u�Մ��\q��8���9��hdkL!�2�j̘�~3x��a%��p�����_��Z#�E�($���܀D�֌�%��j�K���Y��4z#��`��+���la��!~��޸%'|��-h>��|!��3--�<�Q���3��+�v�]�C��#���BH�Q��앱�R�5K�|Ԓ�%�|��+�p_���UR�ռ51��1
.k���p�AIh��Qj���6Y���|��n��B#����xXS�I+�r�� 2�}��s.)���{��<�d)��m��������~����V�ٓ��<i/GLv�P��a���$��[4��t�����,�EgM�i���a{T����X!J֠*wG��Zg�l��e�k��D ���� aT��^�OJ�b6�}nX�z����go�oק��>�>�γ-$����w�r<�n�'sC������׬�_�gB{ݽ�,Α4a��fi�<9J��i�Jó���;X��c�HS8>����B����HJ���<�%ӿO<�zZ,{6٫x�hc�ͧne�u��tvI�,^��0��b��?�'��]�sK��54Gj�G�w�7��ۋ=���y��V�;��1'�� axu��.��p����w�@[�.�C`h�x�ʁ���9ߩ�rt����5�a34H�o�Y��n�����1D����䐑�BD� ٌ]��p]5i*�G��_ih�6��Cp�G1�(d|��>ג�[ɼ_��n����m+�3�,kж���8=����Ԝ:lp���UXB:p�p�ό��Um�e�ɷz��H�uXgf���{i��9ݕtY�'�Z]���S��Q�j4��f�BE��EZ3��1�$p1�R�"c����)�����v�V�7�s��0�,N��&��+
U�Є5~��I���1��\�D=l^]\<��fI�����!�0.�<:<&;��w�,���k_��ԙ�����B���5����u�[5�6�O2鳭%x��O�ޜ,=�^)�l��F@lp����(�t���Q�$	�@:f4E��[��{�z�zv	O��סH�2�z ��
|̪�Ʉ\*�Sv����ĞY���9�Fke���?
�'��M��<Nh���$��g�?7m��3�d['���g��d"m���#�����;���*<:�#��˅b��m�[�@���d�p�1煚&�x	�׹�"��!'��C�9�>?���HjHO^�.��E`Kn����A��]�-�wX�m��ܦ���`�M)"��/����i�Z�2'{�1�^KAM��=�j�:G{;��5��.��~)��a�_V�4�	i�N��{ (?uw��Ox���Ƀ�Ҍ}��Ԕ��2��]ķ ����џʡ)X��0p��q�PW[R�{��Q�Mp��h��R�d�I3�б����<���7�d� G�6hΨ6Nq���L+n;�Y W�c�wr?��:	txy~l��b��r�$�XI
���]��C��!E����:|8���}[���Qf�"���N�G��2�J�-t�IM%z	冽���v�XZ��rE4<W���涂�m��}
3���ya�շ<�y� �J�5�q�Q"EM�(��aE8y��t��J]���4(�1վǺ��3����9�)Y��Y�%ߋx
�&{Ŧ�[%�S���������M��� R��4��r;+������Y6�����4�ۀ���se;�h�`E��'d���e]��!ԛR����_�6]+�F��lFv�~�P��Zܦ���u,�} �p�s�U���
Mn����"� ��ϝ��3��`��㍱1�̕x`��B���#�=�r�d�ɩ�5-�"Ox�tE��9�C��8k�7�).����NZO�1�߼U�c�\];��|l��q�������Xj�H�|��O�F%��X��˹&��}.��A����b#�|���(M��"�N���ڐmͪw�@(�����Ӵ6��sE	��.�,�j�TMd��T�95:k�%/l�3���jM��g	N����#��%���%��ͧ*�+lR[�w��a�ᐱ@�����F�$9'�g�3��7�d_�e�E��s|x��Tt��-y�[rz��]�[N����w������΃��N� >|q��%�MX�%��7J�hѾ���SzF�{t�dpe���/�V�b�U�-��xR6��F��?�EpiE]�n+9Sũ�֏��QQ*xK��/6Jlcu�6{�n�4��/b�#��Yl5~����AR=����z�^�c[���oNjZ��{��M��2�U��w�����y�|K�.�����QW'	�r9Q-�ؔ����Q;�|OƳ�VW=��K��-*(g1�5B�g��9'E�ޟ����������"�[�153��d��'�)��%�U��7���]���:P�岭������Յ7�����E�BԹ!��5>>e�4�|m`��B��C���V�#f�>D"5�Tf3[̱��h�& �5������sD������|w
�Ϡ����q���"��g]�n@u�_FrՑgp�8_�~�Ƚ�{���b��z�G4�)K���<߈FrsӉhܠ����J5����,�\
��'U2�8����Q�81@7S(K�V�zc��ޮ�ϑ<�����*l��(��T]�
byf-��K����M��m�Wl��Lq&�T�1�M�{Rp�?,\NhT�¦�$7^AE�A��h 4�'�SE*��[���a���%/�,%E���ݱ�����;���q�[��X���^���[�������ޝ�������r�Д�R'{9���&:���m����ňo�¦V\]��ʹ�q���g���]�3|��(�ڞO|GK�x�h�?�㹚|01�F��;�f����[2�a[<�$�]b�
J�}4]��8)n�;��&�?%4������;�����}-9[�*��@��s��#rF,�EUs9���޲3�ǩv���.=�G��fs��N�c�/�p��y������bw�O��P.<�'��W�SE�����[p�G�b��z6�j�\l��u�4C�<ֻ�]9/OPV�E`��( ��-��:�45��%�#r#��]jg���}�����+su�������*W�L��8�ʧ�(�1��'h�l���.A��Efi7-�|��������n����N�V4�	��aX
�w!c0�5�u1���m� .}�7S�ڶh{�%��B�?�MO���BϷvq�:>ӥk���}�ﻷ&�Lc̽r:uMއ�ڴ&3f�7}�2k�Pǝp����B�8� UN1ܱ�������\2M�O���ck 
�.%}��fe�
<^Cq�f^�/�+��x���������û����󙨭T^�)�<C��>i��D���%�a:͈*�%�����yTZ:њͬ�u�YT�[y�-W��^�_�����B�%��ߩ5H�Pତyb����ku�L{��u,��[�'����gev@g1��&�L���D�H�%ƃˀ�ʼ��#���a���A'H�8��~P�FBc"�Y�K9P2�&��!�o���Ih�Oe�͇�3C�l��@��BaF�*�=o�*͊�����<�H ъ���/�*暤�>z{�a���u9�wg62�dw<�?Ҋ���#�M�2Z#�$��O�M��CCѠ�?�n9m>��@�;���w��B#�آH�<I+}#05B��4�}������d	s% f��jd%�
G���`E9O8!#籣ɴJ�ۨ�"�n`�
2�;h���}ʽC%�AFW��
���$^c�ᕇ����$$��=%/�=/����s�X��������а �_*��E��o��<��ӣ���U^X�b��7�Dm�K�}�!DX ��$i��U"�p�R<��W��W�:z�iT�3�@���3x�e\���D��J㏆p��^9�L�ڜ�f�/k��>�m�2tB�-��`��7��n�&7��㺷�v�����E��B�c���THp��̥y���@>�@+���v�5*�Z���{�o�����������kc�U�J�C̅=�^&v8o�D{��s�@�nz<��&��,�¼��bR�xbH1! ��m�|���OId�˽�a.8��uO ���cԵX����e����q�m,�6�\�cS�&�h��nWX6t����V��
���)PU�8`�M��+2��)f���Z���m��Ms�µd�J|1`5� #m"���"�!��BH�^���p�L���TTZk��иn�X�Mt�kܑH�V4VP�\�]%�A���hGY-i�c(4�,�$d	y���[�,���Y�{�Z��� 74��}C�!�ޯ�΋��
�ߙ�m�=�?�~�3�]�4�϶� H�<�~���d�&D�k��ќ$�ܜ��_�/ v�������TQ��:��k�0gp~d��:sD��;�2cat�匔챝�)�y��zR@�������q�^�5�4ɞ-�\f�M{�i�A��'!J߫����RX�5�9x�͞<Hۛ$7�M�L�Q2���k�4'��˙J��*O�U�����=�'��˦��gM��T�,⁉����N4�DR�%3gIK}�V��gH	�u��
��0�0��Oz���*Q�~��XMV�K�cڤ��r����D,7�:ږ�Z/_�΀ p����܂����ص߼|
8��)�RO
>��i};�z�:(�Ur	�cHn>o�DM�R�R�����ך�J�'�}T/L�-wY6|L�T���I���8�e�\Q��'���z@�K3h �EE��n� *+B��?�n��s��*�E/�17@���3��8����'�O3�h�z~�s@�U����6�Q���W�p�`��R�O���1���:��7m�ђ���G�Ӳ���Is#�bq�r���rY�U��p������TZ�����	��Г}.������B�\45%dP)A��ˁ�*��
�lf!���,��1\˙l��1ߍ�=�5�B�����eh�T�i��y`��i�h� S�:`��!�C��WY	d�?w����2�dݕ IG\��m[��"�kM����!�����s7�:̙��	�A*���U� �#���-t�.��aN����f�o��M�ji�w.��K�f-�M�i[�0+�e�9 e{?J���D�gB s�]��x�?��ϱJ�;��S
P�#^4="8C���m@�Ǧ:x�e[��F��y�vA��3@/)�\mǳ�hC�l�G�9A�:�1��U�=	}�������B|�J�0c��a�E"j����iO֊a������0.�0Iiڕ�{7d�)y�0���`ePׁ�U���_��:/��l���� 5��z9��_u�a1���]|}�r�:��w���c�o(����(�Z��ר�����w	2��}�:� �?MᎱ�B��h{/���C"�Y�^|�KA>�� ~�I���+k5/atyh�e��T��|X��>�c�pޝY>���U���ٖ������pHJ��C#Ym�/	��D4����Tk�0�B���ihp=e��� �B��5Q�)��&�¸5�K:�p��zf�?9���F�u�
	8�w=!)�?�1+�/�us��8�"n�;�������*�I��f����^��!;��4&,�{�uaforW��O��"�_ۮ�qx�,�}�p`% ��j2�f��[�;��ذ�.wy1��il���101����hXf�H۞u�l-_�]�+��v�E��%~��6�l���q����Ӣu��*�?��N����M��3�Uul_�q��#�x�%�TՉ?FX_s#�&t����}��y8FO���^*��$�:xd�����V��_���Qf`h ͤ�LWZXڒ�]me�n�o�8�<2��RX3�a��{�lg��g�~4\A�ԛx���I���kh�P�?Ѷ"ۻ>MȲ�ۋ�lԱ���6�s5z'Mr��S�ds=�2�9�z0��؍m�$�,ʼ6�ď6� ����Û`mX�@��=�X-�q`ߗu����H�i�(�G�m��v���p��Y-!���(�!�T���Q�������ȓ���A0uz�5��~��p��	-���_d��*hNo�T6��8�E�4ѯRCt,o04&w���Sh�oiI=��Q�f��{���_��6>�n�Ӗb��N�cۢ�7�����ti)ZM�[_�����%����ӂ�@�c�_ӞZ�	s��K�mÙ R�����{���G��˩��?�J���?� ����Hx�J���P��\o����yn��<w̼6��74@����F�F����y�HSp�)����5�i#� �������$����(4,W��QD��gE�L��{�Lh�e�}�fQ�p�k�?�M�-K�W�T���즍$ɨ�`4Z���F��O=����i�h$��{�v~��kt���`nNR�&��g�᭕��X�ư�Z)q}�w(�l~������8�3)C��=�Y��"[$cIx(��w3x}$��'�vG?�ݮ��鎂����O���W�㆕Ō�y��>���P�1lΫ`E��DSg7c��yQw���D�%����6��U-c���Q���)��\�GX ����j�1w�?�#掜���	Ħ%͋���-�Y���mA������8�nT�?6-��DPXWm��Ck�ߟ�z�)�7(|���f���B��� ��#j��B�
ϴ�x�=b~�G�&�� G��[e��#)l�3��K�#��q�D�hJ����#�#m�אd�m�z�F�O��& �Qc�A5&�?�
�f��"v-x0NrV��O�R��A������Ufg�{�D�qp��&|:0��`2��j��U5q�%�l��Z��Da���,��4��)���!Yٱӫz������*BkȦ���W$�;|�(=����XG4�t��ѰJ�#1H��^t�"i�S�k$�{��b�$S��Ѳ���Wx�t���T&e��WX��gOQ����#�����,?�H��
���I���VHu�S�6�69�]��"�NʮK�+�>��5�L��I|@�F�X�"60��,���I�>���?z-<[Q@�Plt���`�jx�W�sI*��g�Ex���Fsۜ��$�k	P 9ɺ���k��H_��k�i�
v���(I���V�~8}$���t4��c��6��]���B��(�ƭ>!��\1� \�(y�GSબ o*��>ē��
i���*����UF-����k���e�𽪳#�k�TCn1|Iu9;���v���xR� O�A~�ڧ/i�'���aVqV+(T�s
M9�Z/��ρ{�`,��#�:��j��&�/Rn��3 �4�Brh�T$W/�I��AiGF�)=u�).q��2r�p�NI������J��H^Jq��ě���TA�E<Za�v&(�\�ӊ��>FU|�v�k��Z���Q�a;�����]h������)}�<�+3�W{z�NLJs	x\A�a��ޣY
�ΰ�\��>l��u��0���,Y��[Z�6�	�^�Q	�"�ƺ*Fe�ʊ� 7�H��k?9�8p�{��>���aL.�b�D">���v��+ 4Ћ��H����m�3�ק�W?���#12 nD��GB���y��v:�o¤�Лux{�|wq&罪�� �ꅐ"�������?�����J��9���Gx8��d��.!FaTĘi�ݚ@��E%xd3�� e�9��;��ve&��-dv$���\�G�_��#��W���2a�k�ԛ��o�ѡ~&	�j�,]��ȸe�[�Ö�����	p\ӛ<�Ӏvw�F��+^�g��M�b��ڡ�o�����s�&��L|݉Bo�>��@pN�[��w���2-|y���i������v�=뵅-���#���sH�s6��"�4��Lٔݎ�w!dg�F3�˟�-5���6��Gf����!ζ
�"R�+�7��Tٿ���<sU��B��C�?��Q���I�ձ7����;�j��uN����}b8siޢS���ץ�3BO.L�3�������üV�jh�I1�@�	%�Ȏ�:oln�4P����	�4\����~�. գ��aw����&�y� ���{�\O���#�
�|[oQ�~���^u9�=7�!�%�8���5�z�h���i@6%���D�w�F��p��q�c�W#��D�ؽd	m�%>�C�Z��oљ�h�����$����̡ fvX�&3ȍ�7c6�[��%e�ip�_�+��(w���H�m��6�'��ٟV>a�K�\��۸d�훾�ۜT,7� J��c1z�|�Z+��oN��sVun��`��<�����	��������g�N�%���F�o!���x(�����!�S��]L�É��.�pҍ�1��g�tJ!��J��{�Ǹ��y�@lcô`���c�_5d��X�F�q1`��v��0�.���`\<1:<���,n�yr�D�B�@\39��� !��]Ϳ���"�x���s.�����T��{�D������]!ǟ)j9�i=�Q
�P�!�Aa���Nɓ5��  (n�w�vH jij*5�G��uG���q�p�����T�+o�n��r��s��.*���K q��[B�թYW�(-eF2���\3�aJ�_��*i7����3��]]�h�q�kѩ��:�s7dZ�i.�s�d��u$��,,zp$�X�L�s}ac*�s��TJ����,�/�À0���`ZJ�]揹�Sbp�.c��Bq+�^��I$��g=�!S��F5��E<�kW�(~���u�,VLȤ��,�M1B���hQ3x��-ɧ��hfˠ`r�xI��+��D
�s���w-�0�8&��K�טO�ړu���9���4X���L|9O�-K���~�op��D.>���.Q�5�"��
\֫uU�`/+�/g�/�5zo�YC9aj���&�T8yϼ,n�}��`7s�FQ���v�s�f�%����*�`8e�k�R���/�!��rN��ߊ�PQEr> ��EPjpQB�Ƿ��3wI�V�B0�����o�#�y��Q��:�nCO�/�P���R�M�w
h��L���N�U��v�Z����ڝ>�:X��<f�7E�V5V��ZL'/���c����<��_���w4��H����d�'Jv��A���mrl����_��Լ�0SӘ\�D�	����FI��'������}Y1��w�rr�c�ڠ@��	6��V�s���L�)/?���2MA�%k1���jc��\�8D
3���ǎ����!��_>��G��.�Bg�h�J�"�R�C�ө�S��p��	�={�H�aYO����v��������/zx�K�:��C�n�}��Ѷwh�c�����^�AP0�Op��G-L%��BN2�r��x�~��&����W�*���ю�?Q�s͙����$|ѺE<�K-r�}��E�O�ز�ɉ{�Mm0p�<s�/��Ԥ	k黂�􊝤wH�4@8�n�|����ɚ@΁$��}�S諣����-�6�`&}�t*"��-@uOp	�ߙ�T��d
i {r�AV�Ҝ�3�'�����=�?���|�j���y�y(��0��F�Pw��2�����~&�p��8M�_(-���8��R@�*�`��2�j�F����2��8�Gk��8eIh�s�BmQ��"��=�I��j�V彖�{�%	NyH7���d�c�%ܶ�ѷ��s�>��E��6�zdD9�.����A�er�N���2����y�<B(W���̽�T�L�qM� �_"U"2��,���*`��֢�'��;f������t"G���y3{�Kk>�nԾ�g�$�-`nO�/��X����Z�kXӓ�2�"1��
�wk	�	oB���<���Ek[�� Њ1�5��`6��q�n�o���A&�"1cDw����o��CR10b�F�"�x�1���y�O�4���S���oq�F�'���;��V�_ ���xj�n��l������l�������iQ��;���jdP�w�{Ȳ�A)|p�
��q�Gss��,K�A�<��lD4���
�aUW(mȦ��H�� xT�����n���x���0:h�C�8����_��Q���_C�4�;���Nu�W_�c෌�{d)�0T���d�#��d���ق?��3�u���/�}�H
}��м�����M���I�6�ʭ�;�-w:������
��fG�X��)c���W'��eR��KR�VУ�ڞ0��S�1o�){#��`$s��^<��=�z 0��{$�#��%�L�J�h1l�jS	�j�x^��X��t56�=�:���j'��K��R��P �%�����u����M��<���Ķ-��
�����@ $�iߺ-*�~��&���8;�
<}۵
Mdz�\����#��\���	KV.�K�6zS�2Ã��?��/`2*/=}?��r��w@9�}T���E��Ue"�ԯO�zfa��y�]8�Lo~J%�RJO�5����<�7W�������P�ç7��U;$�*[�>q.���&�!]��݅>�5�)I���
h��jk
@�x�������L��R�jU�ъ���{���YD�	P��l���r7�&`T.x�@�R����͆�b��8T3m:��m�;���c?-��\ϱ�˿H=�co��f���Tϫ�n���%vL���t	���`܍�BB{���g��D��|�lI�|��(�'�e�C�+0�&K�ճل�7�?^u��R��38�s|��(��:��Dz"niHy�a���C6�w���40'7ԧ�2����A���N�v�A�G��&�,�B��u�ɟ�R'�� VA����I����&��d���'���aѾ�ftM��?���K��.�O
��Qv�\E��oz�O%lw���^%�M��Gw�����6lIEO 
E���9�e�Zk=��ݠn�]~����AGq���(g�%��	����(�]�`������9^A�%�d/S#�����|(�YW��֎����5�n-v�z{:�;qT�uL�t��l�ԇ�j�um� �&g�R�%9(��>gݗ@K������t��X��O�.�7)�e��A��ѥ��#�����ך燒_��}��~��"�.	�q�B�a���Ǘ."��MVT�Au@�����t�2H��� ��t]�h-�>�'���� ��GA����Y䔳��1�a�=�/���R�)�����>�ݨ��+�H���մ���s��P���o��$���8\�6K��9�tVx'�4�ʞ���z|0�K��JuZ��%�s0[�Î�`�0Qy�M�&��F��~�����Ta<���.�Q�<Hs��v8[�S��KM]<h>j���.FH1��Ty��/����˲�p�^L`�z?�"��s�+�����F3^\�뵓�o���0rG��_L#aT-q��#�h%5`i+,�/���V��0��!�ߪކ�<��#&�E� ;V���ܾn ��9�zM�J^�K�f��S2T�g�m�J������m	U��#�$V������m9�.�=h, '�_O S=`��<8�%	L;>����Vo�����p�58T)�@r�<�~7v�����d6.�����P�T�~����8�פ��V��?zA폷	n�*�����/#%[]�,�P��D1Z?��� ��Qب�U�z\�y"S$O�߮�U����E�a��mMȮn8��x�e�MxY��B�YC�I)�η��!L�E��3nt��l�*zO��p˔=��;(M�ҵ��s�wӲD� ��;�NY�&d����U�h1�U&�@���X ����=��n���hI��?��ѕ���oֹ�>?�G8궇�q*�������6�]�D&��Kw�M���EL]���,��`�PЦ}l�����6��1F�����}�'&5��"��dKm�t]���63�8���~+�^|X��u<��@���!�!���^y��D_�U؝�ͣ�6�`ZE���"@�&��8���s�����`'�K�ʉ����xpL���`H|��B����ir-w�2 �O�uTbA�$ �$��x �5��6������q���u�����}��A���S:�k��!��2X�$XP����5gǷ�����*��6�l�1Wo���P�/:�S-�A��ǜ�r���-;t��kfzI(�
W��-9R?�K�@ ���_C��잎�ˠ҇$E�$�������8=����I�A���,�X�����*}���v�B�w��A����뒸�D�v��+��fL2/�B�Y/
�]	�:���(��G)5�g���/��[���y�,ΰy�������l�0�W��oU�`��,��s��*��јBn��m��Ր�#/̮]�=PS`��ٚ�W d�֠K��u�y8Gӗ��o(�b��G������1ֳ����z���>@�� Apθ��b�J�=��t5J�0�7�R��p%ͣ��ʊ�?��	�e1>���w݀��%�Łu����34�?|<��Z�[���F���p�H���g���-��D�g6���}%�<v�Cg(�3ŝ��QABߝ��Xx�W(	��S�!�`������6 �$r�����7/�X`Ȓ.fȔf5������?*d�7��1�wJ�_���:S���هZMs�-w��M�ً�T�`�
~^����ߺ[w�P�W�����M�D1ݧH" }J�p��=l�=�|Qb�Ӭ�b	�Ej��"S;��H@���f;�S�����d�$R0g��%$:���e�W�H^�4�����eģ2v�� ���whR����B7N-AL�	��en_�gf��L�P\��S�f{����Lɧ�k���<��|��,��_�{��(�bW�H�z78��JkdT5h�J�Hf^����_-�ړQ%h��ʲ�i��(�{�pOQ���	��L���=�����]c�T:Q\/�>�����"MH����C�7���/v�Dg��� ��4��r9���c*O��+}����G����<Dg�*?'y ��DTZ%|3��1�-�������	��m�L�qV�7�ُi��p��\����\w�X/8��z�J �)���Shy���,h\�ϗY��ġ]9{R�4�|�2�>�A�@�g2���,�L5C:�|;1��%���7&A��Zʽ��-z��c�a�h+������!��iYK��*`a.��'����>��{�Q�ԓ���I��W����M9���.�Q�զZz<<=�dfX�s��h��+�Z��1��/U��)Rt��)�$�>7MA�рŋ{�ǟ2��y`uR=�\�0��e҈@�n�9v����ҁ�YE���Z)"���"ʮ+I����
�u`��y9A�)&_Ş�e�Y,\�lжo�-@#vY�{&��̺¤ǎ���/�fL͛�c�[���_Qe!,)^�Kƃ�/H�M�yd�ޛ��1�b�������X+E���IM��u�Y���@�a+vơ��/9�
���k�9ԉI^�+���(��pN��t�A���=�[E�S��#QԌ(<����Ï�ei�uV�.	��p�`���61���>���%��n�cR��+��;@|��3��*~�5C�#1J�t؇dZ,����Ƚ�6���Iވ%��OS�:�XY�6�5���h`f���l�2�]�T�4�3��&���!�	�۾"�&�{���ﺑ��>���3�а�oh̢�p8$֔f�G��0GlP�(�4�S���m̈�{N1Ӣ&֐	C�ked����v'�8�Č��ϋ镹d�!���(�	�8��_X�B.V�(}\D�x�� I��m��V�I���UJM۾�WK�vT��[⺗ z�ma���ǁ�&�X�WF��E� ��j 訪�ew/4��6d�Dw1�*#M��+3bN�K��t�������ڨ�w��j{���&�V����lLV�*�8C=�-قg���^��15�o�!<.7����rj�a�Q������t��<��y�煝_��u�A3Hk+���K�}Zm�|x��� �;_ia��;�O��t���$�x#�,�GJ�4G��%Cd�K�d��*�z�(u���*��<�G̀��/<��*t��R����x�L��|��ȑ߭K5��i���_W��w7� �Ů������xV���>�o'�#])d�#?5�ni%D�5>gd�څ�ƿ�7$�
j�jQ̬v\�rx�@aVa7��A_�4%��ĶΎy|��mC�@m��f �P��<7lHq��?��rK~���j?�?A	nH��/0�a%
x��j�i]*��G��W�l����c*"�D��.*�LU�,�c�H�9�é2�*��FQ�h�@F�0/�5�q��I���( ���Nb'���{�8Y�.F��3��8;!+T��R��A0��جjO�*;�aH���^�l��S���Y�[��ܛ�F7�{�RU�Ce���l*�@؂N�y��k>sOx%O7����s����5�Q��?\����@�N>���Ƒ�G���Q�xD�{t=�̗vJ��VQ���q���u��������u�8���OZ����u�.���ؕ���̬Ѣ��9�����k��71��e��B���}!H���x�D��<�i�W.2���A����(�ܕ�� q�C�P����U���*-�P�^�!zLŏ�X�1��ƀ�]AC�5y1�k��I�!qr�7N���I^�!i���P}*J�m��	���H>��#�F�>�A*E�]�թ���Z�
�w�
���ĜU̗��;M!�9�U(k�vjUE'���e�c�vƻ��f�E��1��9w/a�g�D�~��j¨�qsP]¿ec���C��>��� n��h�w?�b�ţ�'j���'��O���o`��KL3^���8RE��H79�fX����NE��x�:�|�5�����\�4�a�o�^:�p?�d���g- 1���G����YO`��'Z�Wi��z3O�36=�J����ÿ��Pc�<R"-�8b\�:/MP:�c�����6�IT$}�cv�@��[��ѐD�^i�u�:<	Un��z�h�O����0E�1��=�vR+Oa�ycF��v�߼���������s~��Q�.w���&�oR��ځ�\<��77���_���y�ͅU~;��S+�r�_U�m���״�J0S���T'�-��
�}\�sTY*%a���9B�Hv�MD}?��f����%n,�~z}�V�O�� >e�)s�Rgڄ��D��w$���́�����L=�3ʂ�EX�Jb\*�����'�A�ۃ��x�kҥD_&�L��e�W�4:}O��6ZV���P��$�:G5[�� �%�"�ʫ���L��2��L&�tq�*?�͙@ק�Ҽ���rn��%��mF�xK�9#�f"zjF�� 	I��}��	���f��h8BΊDK��h���~��gI%�?�w,S�hb�[֌~¿��m�D��hWd~ؐ`�����k��Jnm�>������[O1W��${�x���<̳��F �i3��Ո�Ruwۣ?�|W��?��J������i����L�J<���rj pS� M�^ۯ�&gE����mUת�����i0�(B*�f�����ۆ'%JGꭀs9/�6���)�3,L����L�RWF��~�ۨB�呴�Y�z�?��]2��\b�O��;Rk�QW����t쁉�X�b�����˷��޼gJv7����:�)�5�]��IU�`g�{�FD=��1��Љ�b����x�)�J6M[�&~t)���4/Bf��ẋ�ʓ~�E8���['�yM�ĘB�!N�(agT���	˧��}�$���=�쟺w/�)��6��D�n���@=���L}2��O��Ԅطy�i�	��M�풰q�5,�}Z5�:��z��,��\(�jr8b�hmY�$:%�e*�	�\����l����'����r/�_V�ƷC�O3��ʲ���j+���(���<q��p����v�T�E�ߏ���I���yk'"�G��^zҋh9cB��(U�Lrf[���Mϱ�6���_�iv4Уc:UZN&�W�K5��O��j��ߡQ�՜O�������'�0�5�^"��*W��@0�m �&�c�
̤
ڽ}�x���\�G��'}��YZ���D��C=�Á��;DQ�%�rr��
�W��uy���X�+��F�~ߏ��	=m*����	/_���;U�\�USq`���&a�}3~�H(	�p
�����L0F tdy�<��g|�ޔ��`�./u��n,�pizT�)j8�
D�_��K��ZD�<�o�r,7���?߄^h?�itC��;d���������Z��y?5�=(]�V����e�(R�B۞��KXB���+*�	��%-�yKf��<��6�׆#�f��[��!�x�O�vI߈-W YUV�3��,Ap��+`�my�*2�/�z��C��M�$Z�GC	 ����,�G�
��A����Ai��׼��@e���Gn�M��c{g#b�v�Ӭ5'�C���[y~�߅�����"�<�S7������K7܆xy�m	rsF���_�R@��d&m5r�v5TcN���vZ�Hc��Vtc*������^��7� l�vm�J�lOM��=`c��s����R�f�'���������"�M����,�`���*��+��?+)��̆En�$6
������K�4k�Iw<�Rd�
��&�'4���Ax�sLP(}�63d�p�"�4�4��VָW\�f���:ӾF�l̠R�=�C7�K(Z(��^������S���>ȭ�J^A%�/w�W������xC=À���|a�@u��#D�HCLo��� r�DH|$*ܐ��'�r9m��Q�ۿe\[O^�������	�;�+O3ϗ$��?O'D,z�O)�F�������"zNE������wŶy�_�q��}��v��3T����'��d��D%ܢ��+B�c@dv���+;�q��"�mӚj��c� ��I�ʈ��7ã�&Oq�Y|�-��}U9����x�mFo�q���{�8���`�x���)	�"b#�u�+�8L�$�:ٖ621)�BR�[�8���^貈☣ʼ�屌P�M�kw�Q%���Dg^��#��fGg\ȿWT]�p��m�U�0��/(Vć��-��ǽ�R3ѻ���P¯>��3C���&���p
})�6x$bbY,��i?����@`��,�FVl�H;���E�'��$�T����H�ժ0�h�1k�h���A��^��f;��]Z�k!di=��)���cDqw�@�[h#(�y=�T^e]$���~$�@ܗt<�ě�n�B�~[�ƺ/0��U���%.�Tlw�����8l�ˈ�BB��9���*m�	߂f��~]�$tX����H���ݲ���+�+Lm�w��T&�칙�ڰ��!�Rk̊���`5#�i�����VJ�F��b)cM����7���j&���e�O�&�IQ�d}��#�	�y�`� U0_��hSw;V��Q�n?��ن('�)1�]�X5�k�:Ξ	����2;R���X��J�\�]��Q����<� ��P5,.�D��ϥx�!�ޅ!�� Qv�DZb�Jh�k̈́���9I!HLEA$@�C` ��l��s��N����B`��?z�rw~E��R�����h9M���	�(����OB���NT8<�sP h4v]/�3o�[0��e�Έ:�4�_d�4���p:�'ϳ���9��� ^S�J\�1�:����A�i[zA��:F�p|�]YOO�>�,k^C�w`+6o=�.:b
��?%ʶ75`��������� !��m
��c+�n��g}*	�\��b�"U�뻹�1'�vs&�X �*�(�t�����������¡���BM�h��T��]؈�c��o0	�D\��KaPV��]�Q|����Ai�DseO4�w�C��@8�`���C-�lR���E�	6�P�pP)U�'�87O�S�,ͩ��B����Y��d� LR��gl��j?����giCz F��Id=#��F�ѻ�/��~U���^��l�#39���7Vx�iX}��XF���ڌԶ�ڟI��7�
�~9`�/��7S���v`X��u�Г@}��?��j'��Z��{��l�V�x�
H�ʎK����
ʭ��Ĕ��{O�wv0�U���<l�P����iG.����wԧ�@v�!�P͜U�k�9T�� ���b��/�Z�5����ձӴ���'�&8ʝ�$3:�v��eFKi+�lq-a�����c0!X�e�ڛ���B��+IR�m�e_�S�"������<�Σ0�����׼k�85��ەT�@	�x�^+E�1�ӈ)�ݭO'����ܗ���I��ĳԒaK����vNS���$1\$[�웼f�Ա�1������`���0#ɥ歼Bq*8+��VRf;On}_-�3�xwp�����5Ė��%�n'm����bO���Ǌ��g'��>i�xoA`��D	En=�w�A��c�i�og��wt'"�VV�0�g���v�@�=��k��nB�`�V;e�i�P�b��-QC�m��x-Ɂ'0����G��Y��V+���\�
�z��F��f�;R����@G9�6$��=���鄘�I�1�ۥ�-�A����5�œ�![��/�F���^�W����"�������`��7��*�`aD��t����sI/Q�w��ɠ�2�.��Cga[%�@�)Z�lcyj۠>@6��{����¢t�f��b��$�>6��!nɃ��7p�e�7�ʁ2u����>��G�M-��5��+��T����=�Ӥ~�7�2��꣍��M��ur�E7���ʀu@[3;K�ɒe�vRȆ�tE��n�ڿ������µ@�e){��F!dC.�ϫ%��SOs^�(������/����cx�޿�1/�*�3���]۝���`v	�׿��:K�Wt�ɊQ�쮳~y�o�e�Z:�fت�֎bj@��:�Q�l!���ͦR��X�J������]�<3c|�F�֧�"�Ǔؘ���ُSyR����d(�0���[��6�� �q��%ѹ���V��`6�'��A��(Om�nT�kS�0��\}]�U� ��|��d��M�ca��<�f���B�	�OK�G�o�^��e��s���b�#A��[�\� ����.�Z!��*��&��=��G5�� f�T��R���y�Me^7Ƙ9NT#p��-$,��Ӡ)���(w3�E���U�a�e<TDF��|OIt������K��k��]܉7��+�(0Ii�݇�,��4�r�<
�.)�ʝ����ҹ�_H2\������D�A�#�T�r�Z�l�2�;�����͐�G}Y���oO�V�ө�3�ө$��jMn�D"z�5�Q�m�y�H����Ͽ��j�0߲R�]�+���0��x ���U�I�=Qs�kD���s���L����|����0_E��;Ź���F�r�����N��ɛ��V��/`	������҇�M���	@O�z+�뚛��e��\���8�g�Q�����mq�<�������	N��0B��6��Qo�u�;G���U��� �����_�t�H׉�5З'��� N�@H�J?
_�P43�S��?�W��7����*h���n��I2�Y-��h����L��a���)�b,S��o�8������ȧ���ɔ�g>�������Ule�����"���|��T�c1��<V�!�mB,��{�s���{rnC����s�و��ƕKW��L�M��i��3p/w��,3����@_�^�ˤ!���m��!�X�y�j$Y�����*&P\Ļ�%o�o��m'#������A�=���.E����d�x�4
���*KIz��|a;�����	tL���ڇK���DQ��������t���o0�oS3�RI!�v|Lm�p�8���U-wZ��n�n��
=��B0S����Yo#Bzv
 ��>5|�m+ۥ�����LEW�������X�Z�n:w�Ć�	E&�1#���vuo���to�k9�H);��������6�
%	� 
磤M"e=�d!�a�[��<l�j�&ۣ�'rHG�ipcѸ�P��k�C8!��(Hސ&�`�/��evsq�k�hn�]��R�:��X��<�'O�^�4'5DV�);��մ�q��)T�GD�YH}ʖN�lZ;[0�8wMv&��k����X����x��B�D�5+���`|!Hd��,�)@���6r�ْ�rh�c�"E���7��m�����f_ޘ�:Q��l/o�/��K���q��=|�^@T�f����o[��YY�V�t��>��K���jS�l���.����_��͘�3d%ǋ�l�R����HD�d����-�|�\o���j�!�]�1���{�B6���S�<cͺy�w�^wt-AW׆��6��>�XĴ ��x��ƕƋ��}�f�ԥ\g*����W��1m(���G���3�deٹ���-��[�c��d�7k!11� ]�1��Q�V��03�x�_
�]�5I�/��o���8�u�n!(K�.g�h��?��xq�]m>���8+}^�L\O�IP�*1�9g7|z�h^��[���1��P��E�Q{�;��Q��uY���A��M�fm\�Jp��"��?���/�%�"}��:1�B\+]�2k�YT�4��ﱜ�܍��Mw!�81N7�,�-M�M���m�w9�w�l�b,"6����v��z�d�J-�9��)�9��B����'L�:;q��m�V|;��	��&��
���Y�0Y2�ޝ>��k���t��_SB�s�� 4��>���;\jM��*Zc:�]���-��xiۚ����]at������Gp(�����d)��C�:n�{C�(�tJW�:�*;l�����`�o^�C>Cr�vT�|51���U�,�N֫�(0��
I4;�zg�J�(��j9;��s�fgV:�yF�:#�R��"�{c�aۨ0n�%��C�R@�9+��t!Օf� p$6�C��d-sz�6#֔D���k�8�;oD��|,A{�M�4iK�[���q"�_�vě^��5��'[ӫĜd5VV�p}eoe쓋�ַ����Ī1aΪ%���7>L5,� *)����lD����ǅ�03M$�$G�Dԕ�|Ǜ7$B�
F�q�J���p�w��ˁ�n�?ˋ���`�ԅ΀�Z�LQ7]�l�j���aAq����&���|l���k����?�m�fK��٦]������<@�w�7�I�_�S��w�M�w�Hv^#l� ��W O����ҷ7�h^�����}}���Z�8Ý?�j�^}SS1�P�kJ�rkrں���!�g��z�
*��.<�K�p6W�
��4g���<ʇB���vНHq
ǁϏ=Q~�_F�����"���ݒ%z������S$�,>û�M�4s���5�����3q�t1����_��sW����]|-_0�ri��U����s�*M1��(q�ru�^�^)���n��JCnw-�_k:�g�.�{��\�2�ݖ1�O�	Rg8,j�m�/�19z�t�
�fɈ��V���W.H�b�G�e�cت�G8�C�q�;ʇD� P�H�-�C0��]��f�w�u,YZVJ�hп�.��%�����4h,���ñ��0���N��J�E�m�����C�i�-��`vu���u?W-6v�@��LF9� �����v�Agb
��檆�]�lC�S��Ū�-���	���k��T@�P� rC�+�.��&|a.���^��v^����Hy��CjǼ�ꑢ8:������u��ϼa;�}�k}�_�����n®����G�%vk�v��4a2|�$w�C� ��J'�c��es�(��/����ln'\1IιP��q���y��KF����>V�ꁽl|E�|&�?D �uk^nGm}{t�[yP����5N#^���F/�F�۲C���2�g��@�ԟ(���|�?�y�a��5�7	h,b�ĈBB�������*��L��w�o0 %<�R���)��$�+�K�xM�5f��uBQL�E���C�r
�~�;�猑l�(�L!#�jqr:�����K�^��΂ C��~�=��`�g�=�ބ�qL�:��G}�E�Y�z��PY�Uħ�[c4���Wo^�[V��n��*w�W�I-۲���%?�~�v# ��}O1��� �tNӕ�K���u��Y���k�����G$�p�+� ����Al���q��ߡI��ҭ��^
 �Ơ�*�2X/���yS)DY�����!w�	R�#{BN�S(I�q�^��`ֽ��00�d�=����-��,��"�����Z��^�I
C���U4}\y��{���	���&7�B/�n��5�SԖ�8vw%���w-�rW3pP2�(��b�4�XlUܾc����t��[�&�\���ꊆ@j9�>#X�y�s�e�1���9�L�M���U�F GQ�����f��qH�8�V8�۹L�V����&��U�����5��)B��U�M�3',��E3�x>��@��1�P��r�-Q滗�H�{`�ٖ��:��'�Cy�M���0���]����ְ���.�]� ���	l�
*v\V�I�&x���d�H�gQJax�a ��n�6�ɧ��9����S���.�3^P��O��w�?cr�P����\G}�NC�@���H$V���	�� 5��8X�P�i��y4�r���E���M�/�l��8��a���p����Q����U3�² �1ᝒ��ɸ�G`�*�fS�0�,$�V����}|H�{��Ԗ�9�8�pO�r�;���ݏ���r-*��~q��<�Q�	�\�o
����j�6�|������ʤ^*����,Yn�#ĝ�L��7��f��+�*Rsd����	a�;|���,�L�R��Zϡ��mt��wN9�|5X��D�Z<�i�T�6'c�@I�a�:�fi7㒵��sM�����Ra)�X�s^��Crtzs��A6O?\p���Q[�0��G~�kC���f9>�9�'0M���wt3+�Z�����m������G�D�,����()!F�e��b8�&G��H��7�K1��|���W!��y~ #/��`�X�����K���O^�{�����0%Gs����M3!�tG,��!����*	�i�wgY�QcX��n-sd���x�R��q����۵�b����^���hx��H^)_�>f�?}7���T��������j	&ڦ���_���Rv��Zg�iܖ����L�G�a���{�S�!e���\m�1J�}8i,�7�q�����5wcZU�71���I~1�Ix�W+{�3�#w��bw.�c)1�Q5����l���0��77hC�� �-�p�MK�Ӭp��2���~m2t���s�{	/��,{�e�3 �'���c,��a���<�jɢS^
$*��і�o�0ZQ�����3Ȩ#�+`��M�y/3~U?�"�;��d��q^���i�9D�4�����D��B�\�X�u���ә�'ƴh�����G�Ւ�~�0��L����}T���b�v_��D�Z�8E�¿%��P���^l���B�yX�N�qf���f۩Bc�GXKK�����)c#3�˸u�s�jV�^�(�L�ord�Eu�cA��?z"��&)�zǘ�n�o�%����\T�H��4Z����oW�cj��x��4x#�nb�^7�w�����t�a�{�$b��L���>���N�/Cv'>���)�A��
lf0�q߲ �uO��-O<R��86�Z�T�~h�9#��VK�熃�Lv�S���AXc3Ym|���B� �|�ʧ�̖@��IEvğ=�� @|�g��~o͎E�m�)U��c����ìمm~76N��^TnUC,n�j)�����1wꃋ�S-�j�9�麍3�f���J�9c�����i3
��f�'�du�,JNR���E� OM���� 4ľ/�I;*�+"/B�)����(��,�B��/��5
���l�>j9�qD�C�5���Va�HX���$|�k%��s��+�Z�*Ⱥ��5��((jyq��W�Am2�/��xao��[�s�ɕ���p���0�bH��J�[t��6�n�����`�_�.�.�S��S;��d'ez���a��GZ���'�*�r^�@ף��sb�s��o�8�n�m������x^��E���L���̰*�3�(rv⊰�l��s|�q�<p�0(&A��}�x6muJ3��1 -#��u0r[R�Lߢ&,�܄[�B� �U��>�-IT��i;$
����"�ʟ�_�,���ǘV�ĸ-��Gw9c��D�;��͊5yc~�0��1���*lC��3j��]�>v��r��G��<�p4|��2���g,'V�zj�y�>V�<�%��7��������j��������Cp?�Gr��=]:��	g��&n|u�����f|�I�}�6�9F5�0��i5$��b��i�nT=�tOvԿY���(�L��c.�4H1q"G�:��5 �f��h�LcZL�$]�.Q��8��a:�� G��2��3a���G�[e��0���FH@�`[ K��<���y%�zv�0�wD8|�-fOG9�Z�E�H����. �Av%��q�C�yJ�5M�a5�8KX��q�\i!�XV�փ|���̉7`}c~l����5+���!����^ ��MUZ!��%5��'ͺ�K@�vW�O Ԅ�אV|��!67��o��wR֘���z�&�ޜ�q��'�xm2�sY����dx+��]�(0v"	g�%+�ntB#�Ks��G��p|	0_O"Rl �QK�0E7W��p��;'��2���a�DZDwةu��^v�Q5�?�S�%h�f����(��σ2F���P��՛5_-W/u&�M�����[�^r�l)׸h�c�݅Q�i�ds -�${�&Wk�2 B�Z{����=9�-��Cֹ��|�X@�@?J�ȫ[[�Ԭf}.V-o��V�*"��3�']��a";j�9T�Y��񽦽^� ����|5?���r�B/���&�9�O�͘~��C�.���_���Z@]�`�W=&p��p8'���J��ɩzpj8⚿�[8�������dx6OWrK �����ئ�sr8HTR?��rv/ҭ[*,o4�+�����Τm��B*��%%^ڻ%�츉$)k��P��C�@pW�y�xcZ١B��;����+N.<6twFI�R�V�E{��az+�Z�H�u���T}4�Gq�7���2�n��Q�bM�vb�a�j�tF*��E���8��-���G�Fs�ޡ JLD>�8��e����ұ:w[�y�fū��I�N�a+�]��<���믙�u%`z���
-���1jX7] ��#���qV�+`c$,��1��{��]6�@ *eZ=�DCmMů܁9Hr������kM���0�*C9���!�1ߠ����~RͶvk�.yc#k��i@��Q�.]�z֙S\y��l�|:���'�VRRyZ����*-��6�%��O����Tyӄ/�ۜ-zo��jz�.�m��3[z��?�}C�i�~�_w�v��"�i.2*E�EX��P��\7��G�/ӦҟQ��-��"���ˬ�MҴ���*��A��!���`\Pu�Z��G��8���,�ga{d�FJ�����_���!XO��X��!u��@�A�iK�<_|��.U�ȆFX6���X���\Ȑk>&S��ڌq�)�`/���#d.pß>+��$0��@-bW�?
��©4L8O�t�)���`������Np��͂EZ�#�i�'�i}�sn�! fc�S���/�[% �a�%5�V�Fɻ�c�r`&1*��S�(��r4�����B�I9�
.�A�-�"����3{7�¤��	홅ܶF+	�o���|u��r���M$�=��۪�Q��M]hY?��Ԡk9��x��]=��#(���#Ty�S�
�~��`�#��j�ѥ�}�?8A0U�$2�;���������[#���ɯ��I�C2��#=%�=��'�!��uuBKb�v�s������^�`����&�o,_��Ԑ"mJ#��dR(!2�U���
�p�ju1�C��>Yi[9!�>��>�6���9�v��o���ڮ�W�:�[F+�S�$�L2j�>rT��z:J���T���V��/ґ�6CO�X���<�r��"	��A����& ^ d��kxf/\g/oT���Hˮ,b�:����R�x��,18ǳ,A���L�)���!���fْ�w��y8֟��Ź���C�8!���V!�b�Z�mlyv^fc�rr]\��Ca�ca�8<s4p�ε�q��>����}m��L�!l~'y�Np��\�T�c&)��}d�n�z݂�K�m�H�MDR0@�L!�ĤA�=�A����`�������kh���'� � �}Eg�F:�LTqĲ�b?z�b+�R����X^�
|����������xo���;�WOR
X�\P�S/F%�<�@?�"�PM/(m���O����m
ԡ��;��ބ	G�pdR��L�/�Jz���"k Jp����53�w{]���V��Q�U%�$]��#��`WG�ʩ��*e��ѫQ`X�g�( �.�����;��D����76 �(֋WQ��Xv�|Ĥ[ՃJ1��A)/@=u���i��{�4��^yR�]�Q0���_��Io�l��`����4����������px���P�w���"A����l�,�^Ac�躚F�����i��U�@�jV���?�+�=J0����7��$��n���2,8�\��n���iP�w��@Q�;��OK�Y�a�D��F��V�N�NF.d�l^�Y57��WC:�3��t���G��K��4���+J͟��(����$����
EN�W���ν"-Ep�$r�i��K/�!���<2#I=�u�n���CE�]�M�'|5䉴��Ai;ba�ׄ��;*8x�ڀ����o��ksf@
4j�f����qR�h�t���g��:�z�\�/H?�ޢ��X�垮���!]���W"n���yRa8,�� �yxw_~��J�r��ʊ��rd��t����4V�����p@�1����>�(��"�K���*_�[�H]����gh u�TfOpR.����7�2�����B�,�	6�����	w�.Ҭ��N�0���!ϐ���̽�լO�����i_j[��ʈ��Q�����̔�����U ڹo��V�k�8���N��A�>�ȼ�W�n�t����~��<₝Gs�q���A�;�����kr�_�|��f��OmO]N	���c�F��qàI�<�,�|�u�D�w���1����͸���T�$�#���8��Z4;/<1��ޫ�N^|��t6�ߞ�1��E� ��-
��]�eW�_un:w���`D-���vq1ȕq�g�w�Hݻ�QUg�Ȯ}6DʣR	P��}\Pe�dKϫ�K��eR����M	�dh��/��&��j�t�80&�T Iû���z�!�i��z�u2�>�h��J��dc��b'���k�|��&���_��<p�� Y���'������e�~:ll��>ZPƅz>�)���x��`.�ͯxw�mZ����c(�M��+�Ž�X�C �n����u��+qmh!~Z���KӂƎq��Q�E����&������b��%�X�~�qH�X*��=�}�|*���{{x�@�e��l.'@C����u���6Xܡ��2�X��pOƘ�=��b_��m*�]�v-��IA�]�<ܨ��0�Y	h��~�H��ci*����b�o�e5���m"�����d�Y�"�=퉘�O��EK��5�TT	�kP�z�� `�y�G���i5g�8l�}�C[����,0"��8��7�KpM�sbS����C����0�d�83˲����	�̰K�4N�N��g���Ŧ�cT=�L��禑3S�ag��m^�E.k���͐���ݗ`(�2�Cqu��i-X�3υ&C�F�E��~?{�M�L�Sv�#�x,'Ύܼy��{���`�����p�Y��r'aA�ȓֲ�Oǵ|���# )���S�=;ݎKʚ%�H���x�hu�?� =����	u�x����̳�-/yeJo��ѝ�����aKanY���$�@�-��������c��-N�Ӟ��yj��5��N�P]ll��3b#�l�%E��v�\�n6XkjKBO!���!��H
��K��%������'R��vg��%d�������捳3�ȭ{��/#�����B/���N&��/"�"L��O��e��k	���p*�I�� ?0{I7�TBךfh�!��<gۛ腌���9&`f�"�0;<�_ �����;j��m[�d�pt�x@�-\9���W�`�y��(-Zyz4�O��L ���n�N���u Zu�@dRg�����S�9WJ�$���Q3�-g����qN�ȩ�VG��=df�8]�)� ��M���(�Z�����M~前���Q��,���ю�l���P'�\���T��6[�3���|���7A�$�P�X|Զ���k���C����a�}����G�AF�����~7"��T� ��Qw\������������x��QM��f�	J�G� >��=��"*���/�����t�f�MQP~�7a�`/ԡ�a�C��r��|��u/�Ĩ�#7�� )�Ʈ캛�&�|��(]���ﻥ�^�	�Ծy)�H��'�K)-Y���V��J��9��H�m�4v�6R�:�]nx�I�(�ˆ�;�8�Y�'�o��P�z�z���6�=��1��J�C��/A�{]���$2|��{ ;�Ȃ�f��T�Ɩ�� �5b����5�F8�.c�ta�;�S^�X60�]֌/�|)�;��P�^z�X*׹�3o��'�w:/��{�mm�:��{�f���𠿼�Q3�k"[Z������#m?��8�,�,��w �Ԅ�A��iȐ9����nm2��wM5��ĸ̏�,�$�0p��	�k"j����[������2/����)�Y�;*s�,����ϭG�pO����������̄���龊��A��V�I>�4��T����ĩO.�L��7S�Kr���1�4$�Q�Y�r��S�r8����8+��B�o���+����Kh���b�]�@��	���$�-e6�]t�5��^��L��ܡP�8o%v$����#����g{���Rǜ���	fw�r���z��M�����6����u+�c��io7��$v��#vi��C���I�g��BPK^��1��~�������4r��JPpC���p��_�a����\�f���9eӢ�q��vB�c(t9�g;�R��s��L�]�8��8�Fg�z�p�)�"�O�d�s��=N���n5��� ����~^�P��߉�j�k�*U�}���A�LM��/�IJ�
g%7:1w'I����xw4:����Jꩿ�s�S���W+����hH��x�NXC= !1_�x>�J�%��~�垖E0I�����{`7��|/i_���J��zI � 0+�n���=�tuq͏���ؑ�k��b�K���}Ng�ގ	�ZD��A�8X����o�	%D��R���j!�_�9��n/���N����
|E�<�QϞ��Y���yҲUa���ig��rk�:FZ��̀-0X�n��mQ+=������E�/	�p�{j�P(�0�Гz��&8N���c��2U�{��I��?�#���f/d��z�.S�[��e�-��y>�U�sK������_������� f�C�j����N�k �L��%2�͟�w�X2װ
CQ�
9��U'�j��f���8�w����4��f��%��}hndbiE�CݗI��a���!}=��a����
�+��*�;o�:�2�1&�N���Y��zTG�����H�4xNY�O���K�1�tz�l��(%��I��8��OZ�\�e�����?�i�" �(�P��u�g��@l�T��F�x�V��lfEt����Zq�wu�}ZA]�;y�jWlP�5ڲt���d��ϪV%^o#� NӕG��M���� 4���R��]�}
-ӯe���r���'!�ʈ���.��H1~Q�t��E5k��V��e{�
i�>Ȓ�|C���s�#�{(�a�Ѹ u����@�\� ,vOU���:zO��g ������Ə�����c@#:��G"��W^BWܬLI~_�.R�B��,qV�l��b�RJh�O����,�q�vߋ��5���2f#(>�M�E�9�D���b-y�i�&�ƅ�7�Z���Eno��?�Q��
���5Y���~7�}����_�)$�0<���S����xV3��kE5^�­ə�k��?�bdπ���=��R��|�(s7�a�����Z׋�u&ɢ��Ҳ펥���I	���xH�|韛Z��+`���rX���6�Y7�b�{\����ڬ+\��Gj!U�ʵ���"�׈iJ�ߠe�*��W�::cP���������"�c��q(�=��T2i�EP��;�R�P�g4��0�������vD֟ӟR/F�&t�������8T���F���j���i*�9>�D��|9>��ϼƛ��V��a�V_fO�^n�� �/H0��,	\V�f�;h� ��"�]��\�T��1���@�݌ �7�z�ke���VCC
=?j�v�)Q*�^���Z��z�$X�=-&�ִn�G�Xj)}�&�l�A�ٚ0HpO���j�k�XI6>�	�#���wwku�RӁ'��p���Nχ�+�7�����DM9��,�5�ж�Qָ��N��N��*P�V���? N�2~d�f����eҧ��#_�P~�<�BNq�	� �C�i�ڷޓ��\�$�3����ȟ���d��[I���~R����L��N*���0�%d`Y����7�HGA�Ⱥ���37H�6>	bJ��<�i��Uȯ�>:&q����Z�	w��co�> j0$��ϴ�
��.D��I걶���Wɮ7�3$�>} ,˒pah�@�T�7�9�6I�f���i'��5k��1��*���J��w���̸�L�/��S�q�	�y,�d�.B��6�~?��;�����\*Kzu��*�2�P����#�d�'*�Nz�G��n�&���z����:]]5]G!�����c���W9�X��!D�Y���	�?ujoZ2�Ʋ��<8�MQ-�\ME�x����f��;������t��H"ZH;�w�9��	m�SX�9
���Lc���W(rV0�cN=ܥT�4�%�C�K_�e��K���_+��R]�G�6X|�YeM���T`�_���D��y�τ�< �j�����CI�I*]tԎ�X�hߣ4h�mV]6&R#��H:U� ����dU���^��I������ �[=�A��A��/��YW�f���;��Q5����VO&:�q��f�������1��˜kZ���Lsѭ����Lb5f�fH���Ŧ�\!G��h��	������]���/�ԩ�C
-"b2D�/!]��Ŗ�$��t�sq��\x���K�b�=�~z�y]g5�8��M�Ќ�ĕp�mN������Oy�� �!r5�S��dd�b!Т�_��J��{��l5LU�cw��ZӃQ&r����W&y
�U�g���&FhM���Y�%�J�hkjWՑ�kI��L;l[���޼̄m��x8_Ra|&ǘ[*+t�F1��,B�|�^C~�(Ƿ�sd�eA0B����/ 
#k��(�~��x[�7[t@�}��t3��0���$�E��#ڮr������������qys��ܙ�Z7P�+J�M���>�<�h:u�y�8��v��Yl0��� ����3�4�"��f�"�����MMfm_}�x�lb)j�п��v@�	��0��6~ 1�^E�����#'��t��V�q.�<��?���{��,A�dH;��������,#_�q�y�#+����g���)^SY��X*Zm����g�8e��.�u���1X:b;=�#��b��y`R^P�1�X�z�W��K��TP�(|����@{3% ������2r�qa3&��Q�����碔T�HkM����`�[9��t�S�"���ʧw���B'� �A�z��mG5��|#zl��?j��$WQ$3_�S��3� ٜΦu�^8����߭<�_-o�p��f� 5��V�p7���G.�h��+>
c�'� �D˃�t�X��k��^j�TC�M��L���rg�:Q�\9���t¸%�z4Rht�j��4�C�P"<}8�Ms 
zZ�0������5�����Vr�Ys�[~�u���EGϵ��UU�25�5*<?��C��
����f��Ɍ${0"�@u��.��b9~��ԗ��L#6B\p��s��9�Hr4�C��M38�dUİ��K�ʅ�i����;���l���δ�ؘ�4���Ez4���{�*��A�	m�v^n���P�@�X��L�}�l��}f)���Z�j'�J����?���"����۫\$9�*��I�������]�Gx�[_�2���H�A��	�f�B���`�+�NYV)��D��q���s��fg)(�C5m�"hm����e���x���py��2ڃ����tU��\�uC����\=�d�B��/�M����|aP3l�֪���ïj����t�⫧H�c��f܃h�j�2��tj�3eZouB�Z�<{.����i!�=�ʌ�4/Y�R��KN����q���=����b{����|iq ŭ��忆.K�%�w�����OŶǻ7�~����r\9-+0L�ACmCq>��s�&�k�U��I�n����#����&�n�
�Aϻ ����w�7ut(���X�M ��M{d����O�����Y����tfb ��Z�0�@��嚆vn�����
�Q�����]5^���;�'ʶe���S'V$�|���Ŕ_˱(Q��|K<�B��F^1�?�N��p�� ��ǒ�W�ZѶ��姗sG ���;>��Ϳ����.6�І��n[9G�H�D�30��������z��������vO"�`�6����"�S����`e���{�d=���{Mg�ҁajG*b��5C��Ǘ�ZQ&����Ǡm��4��|�ֈ���.��ϑ�� �ȧY �t+�7E
��?��54(l=��~;7:.Jh#�w�i2��@��2u�c�S�9�S+��m ���#�*�Oew[n"q�Pw�B�JA�@'�Ʀ>�	'������F��a&挼5��j�
�w�V�S�m�T�P:�i9��u{v$?�Fa�9u2V���ph�M�椔�@�W�*#N�OѢ���A���
}w�u��Z�ϕ�}r��=��vM.iI��.���ph>F;����O�Qc�)�4�ߡ�,�[�5T��A�ɢUP�IMB@V�
U1�+B�җđFN6<7����q�_��.h�I~Af�Ƭ�`p�|^6p)�0��X�aė��.�����&������>`��;�$��7����k�7�`BI_r+�1��v~Z�y�,�Q�p{��UyA�!��F��c�Ӎe��]��Ų'��}=C7d�����4r{j�u����»�8�S���Ɣ�|���>E��V)��j�h7��O���Ų�AA�~0m3ʻ�N��yTMaa�/�������/M�VW�����䲡�M=�y��L�H��?��Ԉ#k���6xp�� (=L/f9@��@7gh��]%4iiW�e?�/�.lo��,՗}x� �}�f��B�a^d{�9C���?�Ԕ��f�6ہY\	���
��S[�}�w����]�(�NE�F��-�0��%=�yԄ$��bl�qb�r����"�Ajc-�A�E3���H�݌h؉�fQ���K?�ϵ�����i@4���5��$ 0�HG����J�u��vQ�����A�����rDvG��F���@�ʄs�~��MV`C���_�UO�z�$�w��,���_�e5���@�Ѓq�B�1;'jU:Z{ø')(���у�\?+	�������<Q��������ѝӛR�CF jx_��C׋T�>�Lё��q�)��C �(�8����F��ʤ�%�p�_T�1 )Ṁ�(
����:~y�f?�"F�z�%�v���z�r���G�4�6'�ɂ�Q����ʚ-�@�]�d��m:ו�T·']����0�^�2t,�t���^	1&����J�\����Y`j���g��*��o|�1���G�f��C�풇B�Ѯ�3>�L�X�ݺ��'/#��uIK�Oo��(�T|bs��_)�Kx��0�����޶H�"�>�$�� @���M��s�K�|���O�8Pig2y���'��ŧd�VgS��� *�3/���b�=S�;�z�/,QdF��˪�����1�I�ধ��>_L<,�?���6sBϫ?\���gѺZ
�j����� �=��/��g<j�G��_ '.+S�M��iֶ��וHeu��+=e���� J��.���I>� ?(��PM����^�U�`{�DU9[�W�zU���D�����Wض*O7������|�Ul2�F]C�$�q}�J��.��!k�yƖT��t�.�E."nNb9�g{�}_��L��[R���?ӽg�|(?Q�m6,@|�����C`�R�+�\��p 
mP|���-me�B���q�N�st9�X���ehr�2N���U� �I�~�-�|�����O+��I0��l�5fW����H�g�p��܉\���H0�I�/�m0���T�F�>������$���K���Υ.zB�P�3�Z8ݕj���)+d0�H������!R�+��$��}��$�GB�sr�v��vm͛Y%&I�Hv�}EN��`��Ty�S��ȴ��X2��`!2�������nˆ�eF�wP��v)�Y�//{�@�$ Dmh.�=���>����c4�#�8}��Q�5�_�󜇓�۟≬�����+�8��6Y@��#P�R�P��D@��p����0���?��D�k�=G���~=@����{�s��lND&+UAP�*[���	�m����Ւb;ɭ4Y��X������n�K,g� �C��%l8�H"�-���|2��4݁�P�B��I��#+�U:�+��ز}r���}�Pً�G"�" �m9T��c������p��	񼮡LD�-V�������O3�ʫ|��>|��D4�'[B�u	����3�Xn�����u�@�Y�C`?!u�>����;㋎������{ �܂�n��n���AC+D���W����L J���v?���|�c��yrq \\\����&��9]����{�~�)�kJ��L!8�>��]��^�f�,�LQ�r��f9B�ׅ�+�+��F"5"t]	舒{5�sX�Ř����A�soc�c�y�W���� 	 �����Ԥ^��P��E;�>g亜Q���2P��
����G���^[�����~�/�{�ܰ�s�K+E��a=�����dh���n
ߢ����DP��T�=\ޢ2��AXV�3�H�R�c�a>�FD��S���ӷ[Vy�4��;.Ip�	~�T\,ĘY��tT��gZ�O��J}�wUq�m��p�{��|���0�Y�Ss;�-��
ŉ)� ���:,����D���0�{xD��C�����M1[X��
f�&dh�b���Í3�n`+�A���b@l�xA�^1F��,�o&��?b��� cy#�ݣ3���<��S��p���g5��Q,� ��í�3�(��Ju2?���F.W����
�Z>���O��*��A��^����D����L�DW&c �2Ux��
̗UF�ÿOIJ����G{^���G#!_�o�SB�*Bs7jĮcj!�K`R>r�Ą��A��Ǭ2I��/�Y�:��Lδ�n-��;/�/^oU��)@eSɲ��Cg�o$\�@��=u��W�HZ�C��
Q���ђ-�즲���7�\
mE�t?��m�����0���HD�� ��h��f[�v��M�1�3�s���	�w%&��<�X"��.��mu�ʘ6�a�!���9���5�!���,F��1@��(#���g�PZK2<�հ�z�kB� �/Y=�?�D�ɇS�qf�]�)����}��I��v� ����޲�Z؋��'��'�ΰ�����x�ԕ��n�8��ق���R����&�l]'��<����(Al�jU �h66���Z�khv@7�;%,q�`]��g&-�����y9�.�@1(��2K�*S���U�s��
�z�ƅ�`�P7)z&X[�/|�ק&%*�aN^���2��-�o����+.~M� ��T����3��I�S��\�thʿbI?���=m\أ���%�P�{C���t�H���Z}L�3���]qCd`��4��vS���I�Q��Tm��y�|��A@�����8��k���O�^��,��=��:~3r%��L��ga��0� � o�ST���(�` !��>6)v�:p��+e+�tm:�@��:����!��nRÄ''ӔFyU������3{`$Tf?W�!����3ʊ[,EzZ������,��/,���>A@Q 1Ze�YM�i�Hʄ�IQ��TeSed���x�d�f4K���I�k=:PP�S�^pZ>���b$��*��;�-A�
e�,��d� ��R�%:rKTk�����0�
9�jQ�l-�/�v$4 K�+�BZ��^�Ɲ>品��rE���I3���'�+�>��Q�9�]ǆ�SVpӫ��>���y���P�N��7g�ڐ��@e�����4G�Q�5WJF��[��ۣ�;�� HW�µ�*{m}u����u;�\v���3�L-�]	X�������"jr�+y�I��ŀ$�t6z�l�?��ʈ$�e�����%�)KM���#���@H�������3��0$�$h?/�f�''7���q"7��a�b .��/�����9�0��MN���	h+�T9�1;��y�z�����%(-{Q!�z���y�����J�����.����n�><UhL@?�`�ѭ�٣��ݛ��C%�4V��Ev��ŶS��9h z�����gK��2���O%��ѯ(��0�j�[5����V��4뵏WV�M�^8�oB8"u�a2���U���o�+J\�m�j�fz*q��H�8�-�	RTұhU;���U}=��#�7b���5EʟpXك�����EID2Ѻ%�7!����5���_���:�τ�4o�R[���Bπ1(�Yn�)�� �H
�����xZ��B�%��/�SR�=�B�C\t�i��,����U?����� -�`@�$2�Ӄ��.��2-ʃnʏ�ls���J����8�_$������[)���UL"�'�Rn}�m!U��Ν�kϔnO���H�NPd�07�*����K#�m�� !x _Z[7���.�0�R)��@A�y|.��G�(_݊���8rv[���N�����;fB�(���*��*��#�������snZ1~7�I��}|��~&��Mϯ `�5�% ���^s����g��8j�N���/ �75���gF���nd�G��B�� ���F��D+j�,��<�
vcг�=���{�u�CK�ցD�x�Y����prV�}�t�f}#�.C�W%�Q�n�QJm�U�'��Z4���mMT����BP{ڦ��nz�H)͆D�y��I^XP9u�B�w�W�s��Foz�͙�t�m���z��'
$OjRU��2A��aJkEn�&�����3�:*�}�yL	����e�=t,���w|{�ax��BO��&�b^����8E�J����������6�/-��27���g�R�� ��72H��C�4wm
�0[J\�f0�.
T!���?*ы�9965�l�P�'����H=^�0���?�0�2D+i���!=�8VX�}S %�q8.�`��0k~?֊��Щ�IJ>��m����N�t0_R�67�����F���|�����sd�G馎����>R�aԀ@H��+�w���Ѕ�3Zgv~�{�&�s%I��ۑ1��0�\����_�:�-�K��p���/5�4��:��o3�fImy���c��m�����[����g7�&�.ص���?z��4��c
��Z�z���U:̀�z�Z)GV�`�>�>����t��xG�c�����n�H�F�)I9U�@���gk��XuΘs���U?�j8ՠ���^���/����k�;4lLe�FV����(F�Β��cz�sޭ���YAV�A�)P������1����x^���+[�.��	i§�fξ��`	��Y��>��`�Y��N������a}y�M`΂
8��+t���&�4G��7�^�Z����d
1,,��w��f=p	�Q�%���0	o]��a�R�'�_r������V�jb.N�'�=��~s��_(�[`��K�͌�BN����!��L�ך�QD�c�B��Y@��X�CvoYsW�2)��3��F;�KD�$q�<��i���M�6x? KS�{ �,!�e�=��_��S3V����J�쬛Q���b��G(A���n����G�ײQ�Dy�\�F��a��7���ѡqg��fX7�,��H'q��q>��{��&����*|�퇂����_�(�AB���tF�U�T+&8�?�����Z��!�D�o��+
ס �;_���?�4ڶ������Zcp�[�F�q_�Vŷ��ȵA���}�*m��>�B��[�t}hڈ�l����]�ꝮI�x|�cȏ6����s9�l`�Qw�/�D�w}?����r�i9�H�l�� H�Y*,hr�t�|B��3��^������"���.j{���V��wy㥈��W�'/�����M�(xП�z�P�M�k{!`}�?C|�?�Q��I���GX�1��Ɩ'������j�!G�����l++ECX�C��B5��=B����ʍ{���S>"�R06Ič@�^^��z���Hu>�x�CJ������4��J��J+'�O�;�*��F6jCp��0m8��藞�X�FNI����hM�p���P�	��i�]���3�9���`L:�Od�dKb�>���s���m�2'����h�2,S�j�t���s\�>���=]��}���l�9-�0�X�`Ů���Ҝ9��r3��m��<Ƴ��٧}�@kFl W������ذ�mTv��z�ý�>jI�=ٕ\ІL��a� N��-y���?�4/�خ:B+�fm�������I;.�Xz�t3~K:�[��/�s7V\8�$*�G܎xH
lz�&����64�°�����Q:*�
Y��A�[�z�Ɲ��N��攣rrC2��z5҂QD�,��PY�����	�*��t�^l/���)=Lc���H"]F��5��3q�H���ơb�Z�����[o�Y��dNa]i�@x��L�ev2�f�a\|^��x���ߑ =FH��A0?�ח5M��C�4�Q����P�N`�=�J��u�i5#L�P"Ls;�Κ�Y��ku"��R������1{ۣ��l��}��FMն9Q� K�j�Hajޞi,.Nv�A5�.v��r��^�W�b  ��>�B7�60�"qw�����Ŕ�ū�636�[�	}��>4Y�r5K�+0e4��8���`�9)mO7�Q����1(���U(Fe�y��B>�3�C�ҒF}7�̽[\�@VV���z�viD}Ym�v�ܙΡ��������%��J�G�3"�{7vH:���/�c:�>RR�x-GЕg�����emƹpA�,a��f�b�졝�Y���rF��uޱ��hG4�
=����೮X�_X�s%�Ch�މ̞�r�Q1�zu���R�H�~�{s��m,#����� <X'=��'�Ƃ =��j�&�-���%ngL��l�qTzF?*�?c>��v�}2"O�:Q����w���~z`3
������P6M�"��&6�l�<�d���
}Ϸ(>�^��u�T!=ek��G�!)a�{F�ΑWŹ��
��e���W��������T��]^}�5N����~^��R�Q�%� �|��jxW0����A�>����}��чCL��J6w�E=����[ut�Ȏ'Ig��ggɪ��FeƦ��,�zH�[L��Lw�Jr�r"0��FƳ�!lQq���gZ#%T��9�BL���@�'�f�R�H�!w#��me��eE7�f���]�\|T���xIy��W��wU4�^NH�,G-�erA�̂J���ڀ���U�}��m�t��*�j�Q�)�L�'��0��w5;Dʖ�ϗ��b^Wz���B�q1�\/|z���\:�cݽ����<ѱ�����	o�ɜ��0Oe90�fA%:��@5B�
F�{sבI<�9Zk�a@6�P��@���DR�h�z�'����r��[� ���I8D�9v�L���"�)����|D��0��_���&�+�f��u��B��s�E��G)���!��xdٺkNbY&=/���̯���5W�����ص{ٖN��;����L>��L#Z}|@e7����%�^Kң^�ss�@�X�X���(=w9NY��m\����-�8]��VH�=*�G^P��b���9L����I]�62�үa�ĭ��Q^>#��qI���$�n`�4PS�7$��C2��S��o�R5��}s��ϒ`\L��h�[<��{<��'��=�#/��
߱΍=��Ʋ��T��J��'/.��`�@:/먾�m�g6 můq��<ڄ=���R�{MI#���i�05����D[�*�{&{v���">�w��2���rU��g\�x)+t��� �%V4�%H�Fѱ���v��ˡQ������Q�/�y�%h��.m ��EP&��T[C��HO�y��U?�����4G��h3/�UW�g�X%���A'qZ1��>�F]����hȌs�S��Xǩ/_�k� 9M,���f�#Vcms��W�a'�%�(��[R��%{@�h�����OuF���j����L}ìJ\C��d�4�43�|�n�H���g����b����U��O�-�����֐��{�W0�ى%xq��e����:кw�yzZS�i��]��Ͱ�T�<&���
�Lu�-��&�M�n���r����T�JT��ü0�O�xw��Ώ�1w�?{鼊0ذG�?L��<���!c�]ˠ�����=�-���d�����+��U����8�DV�ߥ`��9�RS���_la���\}�%S�2O��B�=I�C�UԍdҦ�'��Qf�F��CK���ډڀ�~mH%vs�q�1p<Dk�趉�F�w9H��������*�"��L�$ &f�72L�-�ܶ)p�E������`q���郛`�)V��a���ˤ��h�:K5I�[QoM��3�8�y������D���(��{*�mo�=^�܆b�Co�tk6����c�45��>0�B��5��++�c�ġ����K.�Q+�H�F%���d��`͸j�˨��f�)+�\N����w\�(�su�������_� ,�UD7S�҂;�%R.��hw`wy�qY���X��n���(�<�����(]=8���kF#�Q�
��9����
'x�/)8��4��4zP�*���H��_Nj��ܧ! -�i���w6 ���_a�`�!~4�D�ZI�yfz�%Z�֘�e��}g��a-�t
Q����*��(�Uu��ġ�)��V7C�{��2������_4d��:P[*��$��V3��s��KE:�RQB�5��� !�f�빽�wfCc,ZM�R���-��j����e4���9�p<��Ě�U�/���Vrj\���ރ�&�Z,͚q���*��ۀ�J"c����o�!��I;�4��XG�}d�Ã�5x�z$.6ȝ�`H��*���j�J�����B�c��"��R��h���ۮ*������Q>�^7�6�)���?��
~�f���Q�վ�VT��n�鏔��J��K�i������=����֓7�p�d���#�a�:.�/0Ldx�n	�P�h��Ǆ�l��~�w}҅\��R.����d�_�5����~�n�)b��Єt�C��m��2.������YBjD�c�h�2>S{#P�C���L����lB���*�'���4� ؾ��w�ҹ�����z�dI�X�����\���]:Ŝ�9 �/�Oao���Z�r���<��gH8���l�K��3H��_���	����]��A�2��q�	)B�>��鮍��A�,u�}y#uܞ}�����,�bU���j�
hn䬎:$NE�~�u��k����PɅ���z��8/�l��a�Gw�ؓ�)��������!Z7��c��.2���]�����(6A+Z��S��¾l�F����-,��4�����Ѯ�wR=ˈݐ1�Ba(�jK�K��A�!����WM�ڱ�����&7������j��?�T���JF͙㿒���~BZL"�u��n��.�j��B񅽓@]�~�V��1^ٟ���|��6q��F;����pq㦷��l�l�Jڕs|?.�5�|��]�;џ��m���͖�ت�P��p�}���-x��rЯd�y<�A~߬~3�So�v`��y1�æ�F&'�z�-R��_-��q�f5k�할�*b|��q5�3����&v���*�nT���{;��.���LUܔ~>���((�R{�kɇ╵Z�������~��]:������6"Ȕ��a�KSq�"C�M�ma�0�A����m��~'��X^�C��[��:��e�4���07j�o���	9n�x"@g$��|��6�GF�f�b ���UlSr�������\��M�$)��長4z(����U^.�ƽ�'\{;쨙�c��",���wtB�4�q�if^�6��1hd��2~�q��+D
�1�I�j<�<*cL���U���X���l$��\(D
��m����Civ�I6��Ԑ�k�8!p>�=��?cH8���Z٬#�X?��H�^�]n�f�����83�M�����b�P%K�F�H{����s�.e�K(!)��A�jV���X�r�i��I�m�Y����t�D���Q�#n���6��*��@!�hqT�V��O7m���M,�&s��q�ݿOhV��»�w�θ:�Us�8�����V���&�K�|�C&m&�}��������^*�SyM}� �x*��n5jY��(���ru�����Ǵ��\X��ǻ���t�Z����u��0qkF�˦�/֟�6)��u�&ϺH�
́����E�nn�/���	���#0�}Їp^�#�7F�h��K��)�γri�^G�S0���b�Ȓ�t�d+�?����ႀV9�� J�aw�����Mэr$�z�g���Y�%�օ�E8$�`Uq��~�;���ڠ��h��<8Au�*l#�T-���_/���=�[�fr����S�a����C���o��JQ��>�M�Y�%���W"��V���G'i��Jg�&���A(���]����+�Y{@�ښ�c���JYƏ��$;N�Ā*����.o�(�������(���ܲu��~���_��SH5��T,\}A�@�K�) ��*�O(�Ƈ�_b����m�j$۫�hg� �?6L��J�vK?�����z?�>�@Bc����߰#�|.Q#�ԝX��,h����w�4Y����ձ}��rW�L@��dS�+�7�j�X�*\@7�p�}�Gɩi}�.N�����+ű6��z1�(���EK��*��SL�$`d�s��Da�BvH���G���JW� �7���9b)��H��1�"q:����EB1��orc�Q�&����xh�xtEM�Fׅv{�C�f�C吤�N�k;p�*�?�`�w0�����Cx4�~�*F�˂i |�Cg:nmD㵎�Ƿӑi�0�D��i�|��1���>�C{Ol�#b���JB����m)��ٸ]�7��W�\#7�0cN%Y���lY�d��!���:�˲I����F�:|�$����Q�Z�~!������Q�"�(Z�|9������t�@xԂ�/=uo�l���?u|/^J+Ih��Mf���O��f���|���p��Z/?�}ldW��T���IR|ڝ�tl���=�Aئy���A 	�H`��[Мܦ/�j_�� x�2��s% A\��G|�������,���*�~x�/*�!� �b�Re�̊�JH�4
�Kp>��89H�ϖ�t��ߕ��Xm#)i�	�u����v��oR���l{XU{�=H������ڰq�&�	���yטQXP���mr��C��:zg��8��
6@P6>�O�E!��Op�cɢJ���&��b��؎�7����KO5�@͠+�iu�wx@:?Q���.p�閽��,�@��q��j�z�B���[��]�^�zbX�SJ;�7sg�F����ܓl�s����������r�����7�-)
v�����8�(�
���;- Y�5����Ԃ��³d���������	��Wح�AI��M4��ď�
��Ѳ�Q�SWQ��4��*��@��,G�h�Gr�.x��)_��lC꽿��S��:�q�+�'OrH{'�>�˼�_��)�,Ō*<�g�
�K��.8E&3?��dp��	"�Wt�����w�����<�<�����7 ¤U�
g�+���D#�X�VC:��.L��L��[9.PM�J�	c�F�	�V�3�Bs����*a��ea�j7���>|V���ʖ�
�HH��"�A��ͅ�~C~r��628����Ɂ�T�(�9��D��ؓ'�����Bo�(�o��x|��T�֩�$`c�������eҶ�f�@��%�U��}�,�d�*/�a�e�2��tta�5*n���G��\Ҙ��������I��Ol}�L�a�@�#���|l̰O�S��-�7�X<	��o�&`�#�C~�T���N!���3�~7�	շ���קwÛ�-Rg!f�6�����h���Ïh�j�����h� �x�ʉ��[F�?7�ů�f�	��m}�0y|ŧV����PY�D���$]�ld��$3����ldEV�	<��	L�6`����������8�u4�:x`ﴩ�ݠ�
�=���r�;�����Q�̜6�����aC-�2=޷��=.RW<�h�L��A'��\��)��1��2m����ɐ�*��3`�R+�_��fn]L�c�&~���3r)v`0e\�gBm� ���g�Gf����'O���;�T	��*m��ט cp~�O<�-P"�n�[v��]��ޓ���|�Y��ӱ;��!qm�"��D�3m0b��Խ� p+�Ģ��	F��-S-e��Uූv�Һv��ߣ���F��xIw-x91�켖͉��}9ʩp�ѿ�Ϸ^�=(��J������h�$���[�A ���^�'3�1?W!sP�c��.�A1�A�ZX�L���x�wn�@����
p��4M(�q�d5wb��k�-;�h������X���N�Lx$"�\e�,}9�����.�ٴ�;���WYYǳJ_�;��1_��e$��l�DQ����	f  ����*�&�:E�C[����_�/��0�gz/h��|_)P|!�s�"��ʑ��hiͭ�2�c�I���^j�_A!Q�='�^������}΃Px�FI����э�WL?�׭@<�؝�&ˬ7��[R�#�VL�Z�m�{�O���Ə���l�
�6��=3$e}��_����mH��Yn���ؗlCi�L"֘b���xj��{�k5����B���u$�)�&&�G[Z�4���R�y(!H�@�~�@6c�WD{��OK��D�&Jڞ|����\��o���Y,�+=���ɂ��&�(��?��D�ɽ��Te`x��C�_�K5�C����$�����Y=�R�L���)Kq�i�m5ARѬ�0j�B�_�۰]�n���z-�����vm�a�����@�p��%�s��;>�x���!��z�N?��xϴ���'֓����O(�g��||w��FW:���a��A��Ϊ�O�`�ig�??5D!7���%N��m�>��Ҹ ��RY���#�<�0`(��{�||,!��O��($ʆ��]ӳ}�M����=@�E^U�A]#�9�Xij0�A�ٳ�j��ϸ\Ŗ�+���cN �}���y9f�仰�����y���Ui��R����@f��,N�ᗪ2����>!"�3(��i^�ѫu"b��P}�+�����.�`������f���+$ޡ��������P!��U>j,�����]� ¨9q6��ʅ��g��L�,|�c7F}=���`�a.�����F�o"��N@�޵T�Rg���E�@t�R�K���Or����϶>��UA���
�����)/�]�;���m<j�s[r
{
��>Ƴ�?ŭD���m	��,Gay/Lc&�C�J�G;R,��L�QXA�����m����C&�����m#d"��'��@��ѵF��4��r�%t�����t=��_%�A�RW���EC�ِ��ƣL�oЛj�G_js�A	�-^�gW���IrW=�*NƊHgw	�W�U�����f�"g��r����XhڨN��buh6� �VH�*�py��f���3fx%�Cl���_�����L��A��u�H��CjA�%���.^�l������7��J�F_��$
�e��=�lw��PLo^q��Ҋ�×�T��F�1���V;?+�P�B���*�����n����I�,�v��8R�w�E#�����8>b;*w�E�S���*7�|
��F��A��+��j��'�k{���=+p<g����7��&چ���Dp6f��3481�߮m������J����sց_�pNY�=������X|���Pj�mpS��N�l�ڥ���CH�!�!�]i6��rܙ��z:���@���健��KmqH��d*�kR@34s�[F�в�R�E�x"uo�&��Aء�ʛ���D�W�Gk��S#b=����T��Y�6�vV�T����R "���ք��f�͵+w=����eo����;�l�\3��%{�z��$BH��2u��Z����Iפ*�����j� X��R&z��	�oN;���1霕��E�n���6�~%���[��/�"?���/^rP��V򴊌U��3T��������7^D�e�IMA��P�Fj��z9��Pco��<�&����$O+�B���;�l��1Ł�VV��r����.��	� �h�u��'��q���z�s�ف���J.��bð��~A�ۨ���s�YI@�c������$�,�:ی�?`�-2?k@��w5�C���R�Ԣ76�-
��ѱĉ�&�u���I�_�D���q{�*HGw��.|ɘ�Z�I�op�r¬��2?'I��A�;�mi-��+�"���VE+f�lZFZ�a&���S�6�e�A���Ǳ�\��º[�O۾�Q���.$�f�t,��h�������;�����Ј�VP1��Su��&�M[��f�X��j�Bj�T����,��\Diq�c~Bj�J�����*����hq�A�]� w�i(T�� �_��
�����8�e�J����$˒E�@�,�U�)��5��;/횏!n�L�R,D=d�^�S+{�"8�-�Lk*������Ђ%�_��^���������Xb�
W%`��F*�6��Qs�25���q�p���Ɍ���K�j�Q����n� ����`RH�'g ZN����j�~)�	НWx�6D������2��<�x��N�/����r����ԫ���u���[��},�S�멝�����O��R�X8�"�v�No���o���^W�v� ���x��u�A/�G97��2�\@�A4 9꫈U�0=��U�W��K�p����ɲoyS���,���4�o����=�<X�%f՞1=��ZВCnh(chf�dw��O�޸�LVO�SA�Oy˜�:&0߈n�>�<7G��SCn��*�z7��-H��Ԁ)zK4��-�ʎ�쬮��b�A��څg��vJ��t+��賚hӧ���
n�~��Q[^}ӻ�|�JΛ+%�x�f:����V���أ���6��i��p�a��j
��os���I�ć��";�u%���?�v��p����Ć�c�d���`�B��$��������1�q;�`��>|�dX$:)�4O��"��Ҏ�j,���$�*�5򅎸�.qRV��O�l�;�x�0�/V� �A�1v��-�wIx�ɝN[䓡ńr�D��O	%~lo=|�{�R�"뮼���#k�M�/���Bp@KӬW�4-v*Wnh'>G樶����L�S���������c�Q-U�P���R&`�E�<B8Љ3���?�̃�i��s~�Q�����-�J��)��xc+�jvDp-�P>��>g2N�t�R�*Ҧ\�Ȼ����5)՞����QH�(%F�H�H�����pC"<+&:�O)���AKoA��7XV���"^��:%��	9��F��p�,�������
#�Y"g	��_�%�J:c����:����:Yr�_��)O-E'q�:�L��j��z��?�a�bw�<O�L��?�v��t�&�t`��_�rvN�RM����Z�e�"��7+ಸ$����9�r{.K�tn�8ɩۛti)aʗd��_���TVqڪ�V�o]������\>�p�s�c�	;�T��~a+����๒��O�A�z]�o닷�m���G_���8A�l�
�_����T�^=E�i���=&��̨�Z#���K��#Α��f.=�����e%~��Dk]B�1Ba�\u���<*���7�����A�5��ƷK)����Z��b(� /zA)�x~�����_g�;Wz�� À�y͊��AQ�:��q�Z��z����%Z
ވ����vA�����MӰ�G�g����Z`��F�i�����96�克��WdI8�ݱ|И�u3�ze}`����� l'TZ�-��jϴ��<�n(��7�o�:5ޔ������<�ʝKSF�H�c�U>�+1/$H�X^:v���0���$*����ЫZ��	�fob�/]�쉷���*8_@-�k�U$���}h�[?�\{�C3�UzN#��[�O���5x�vA��g�[S˰��=��n��h!_��
0�N�O�2��d:ۏ�H2h�����+j&�~��/�C�����g�٫sY�OE{u��DK}��~�
����yI{�ݣ�S#{p$�z��󄔱�&4a��=9��3�N!wS�g���b��IP�~���b��P�?d����Z��;��j�WJ�pL��r�v��Ğ��{�Ų9�P#wJ�Q�W6�iʑ�	�W���B�J���z����p:�K��P��=6A�[��MIJn��ؓ���x��=�Fz�i}R�z}m^���cv$=�<��9���1�]���տ�m�9�����]��5j"^���]�j̈́o=�T�m�����XX�ȅyi!I�iz.D���S���S?�&z�ܑ������]NQ��&dP.+��Nגǀ8ʸ�&��N՟^@V;��5�7�KmG͇��0��!<�5�@��"%1a!���J��E��",�J��zӵ
�'B(��.6`�u	�]$r����3}s'�>���U�쯁I�Rwm��~��^�{��;5������OJ(�:�A��$v�sj��F�p����b�6����Sڕ���U�3ȟ����ة�џ�*@�E������hnh@3�6<�T��${K���C�G^D�Z���|���Wyܪ%
gv�l<;�K�����C����3���'h�P?[�''
3���(�*Uy讛S�Mj7�-�nu-;���b$|`aǱ(ؔ ׁ"���nJS��5|UœEy�kʦKN0��YDx��N�=T�NP�9�M����k��ޮ�pc-�����d�(V\=F
a5�����5�v��R��C��e� �g�Z2I,4Dn���H���E(w����;;,����1��c�	�<�^Ġ��9��\�����[á���W�TH��{r�����O*H5
�=�!^j����6�!��9傌�g�~�<���[_���8���DB���+w�3=��h^R� �Q���a����B�G�7Uo�:��m�f�咥��fӤΕb.I�2���S�D��W =����Ť����E~̈K˕�V#x�R��Y8c��(��,��O���Z{��ZЅ�djk����l�Q�Z��d�e��������-�|d"?z����?a�n�Yp�V��B<?�����ɯ��o��Pu�I��bά)�^Dٻa0ã�/�GXu��x�&嬇קo�a!�(,���� /b�/�V�y]*~��?N� �P�gGI�*���x����KY�-�k� I��G8\`���Յ F�������l�uQ�|�]J�\Z0��I��Z���<���
�����F��\����v�l���l$R!ֶs.5��!䟗���fe�p/����HNE��0~��UE:�^��B��j�)5�nx7�M�����l0���E;�w����IH�i���)��e�>����\�u	׊�3͉Ղ�J�p��s���ܳ�֤U����q�ok��=�E('��HRV�渻/��o*Q�+~猴X'�_I���]�3����(:"��$��i�5Ѯ�:�:�ll�Q�����������a�&�����S��ވ�z+�8q��V0�^8��/5ە(��v}V�l¬�W���lJ284=���tA6�h�Z�"6A�=�����n� �<w��,T��Y]e������8)��Z�	���Ճ�\��%�� &��H���s���Ī$��.?\�F���l�'2����KQ2wGQ���i�%�LEW��U'����x4j4��}��+V����������{�hG�2�K�d�%PE����
�H�G:�_b����qJO6��9��rL��M�����;St�z\{xF��u�5XIO���JWP�&�d|`�T�����R���&-}�M�"]q��V_˃�̱N@ (�Lc��_|���T+�� M`� ԤVZ/��ކ���8�@P-Ј\����RJ5�3:{�C�x�����eb�P��xU�F�w-C�aB�A���������#�������.��#bc��4��8A��G��B��+��R	���wKv#�V�D`qc�c?1R�V�mﮂ��5���/�g���9_{�&�3+7%���YFh>:X��j�S�K�q}�5�/��Ǌ��&tg�����=
����)��j&�+R���&
�_lI�bF �5H�Q$䶫������C���d"��it9UE�BT)u��@��4���ڜ�Mcߚ�3���ڔp:tE���S�7�VH���P�mk	^�m��[�}���;%���Tc�nlQ� ���/*s�� ��v����/�Ɵ��uݶ�G���s�i�ϖ�uGl+��=��WT�Ha#4����u�Rߒ�D�����%�D��Q�g��h�Bo��}�r���J�q��އ}7�^�̅J�A���s�6��Ԃi:Ѳ�ۢDN���$g��}ZY��PtT�^���ە�9Fn�e�5���A_t	|��k .�w}�"����S���`�E�n8�Sk婽վ-�=�?U(����zK �ٞ���E������5 �^d��69;W����xF��~ܵ�Q�{�/Ɯk�<��@��'D�,�L{@�� ��?L)�@�sO����|�t�m[O8�!�Q��l��F}H_]����y�e�zZ�Q��v_"�u��g���#�G�q����r�yr�=ϝ����T����S�k#��+�("�dQE�R�C�b3ǻ�@�^�8��C���7�6��YKp�D˪D��H��Z? ]Un�#�o*������;�ځ��;��U�ԛļ\���*2l8<���[��K�~n���hĠZ���5���� r�:��zү�P�A��8LE��E�I��d'�y..6c��p��y�E@���Z��7�6�'x�uW��/R�w�d���*�z-��g6���,{8�(%!��-e�9�DZ����h����Wﹱu0��R;[,��*O+W[�w`#��U\r��u
ۂX��Ě�B�υ���@��b�8~Y��B>v@
HCK��3��S�X�|2_P�I�� �����J���Gi�,���E��]=T�����ᢥ!�Q#�\� �ú3��6,�^�����b�:��� ��CƩ7\�U
~6������:���7^T\�{��k��0fB�8�:h���t���[�x��e#��� ��^�9U�L����m&}�K���q�G��%6�������.���^�<ʗ̂���( l�g�3��]�B�9��K�s�T.E �+i�9��ۀ+)��-���Y��8x�,Qp6���/�}��?�s�gݩ6�bV�o�~�G���>�nS5��,_�h.RUk���Ꙡ(��B���x���6!%�e���$���$��l�[8���@Ŀ�����A��x� o���d��}��7X`�fM�ތv��l�?wkIA���T2	�t��vaɲ����1b����T^hЂ�R8�5�����w�pV��V��a
w<E4�P+^����pA�DEr�[K� �l�#@=:���b����]e,�Ɗs�Լ+g"_,�d��m��,d[X�(!2�א+k9uځV�����;Q�E�n�j�u?�t%�xQ/=�3n�<��o�{�
=��|�]�U�1�����x؇xj�=I�rQ�u<��vy�Y��M`�l���F�c.��n���E�M�¡�.?�J�v���̍�A���f�'G�񀤫"���%=�nω�u�C����P�ǜFѨ\�������<��)�1EK`���Z�;(a�P�l%�B� �;�^^�-�o�5Y�i\�ir�c�kA�[MEJ�d�����FRt�ۙ���X��fk\5�v��{�Yc�!/�cO����L�0a��e�K�9����M\5�7�&�O�NKx���k=pI5�Ͷ\�ݷ��J�o�Rc���<���٣�y�ϝ�)Wͨ��I�3Zi�.��;�`L���\�=�]��|���
����j��~-��&m�J��fC�6����%���6 Kx�m	uu�ؘ�W,�4��)S=e*_G��)� �z_�J��|.GxeT@q$�_=�CU��"�=5�]|@�N��v�W��"Z�+i�׻Eճ@!N�vh�Uޟ�+ƨ� ������jHC�h��5u5���2.`OdFAW��XkT�J_������
��	獟�YS<�t�z�u�Y�c�ہpإ ���kx�����!EW\^��=��
3��Ӛx])��Ғ�$hs6&���o�3�5,��.�=����T
������ ��}L��Fa��육^���db�#�p���~���S�
�;p9bR.X�Ŭ� %�l?��W�3@�6x����tv��B	1�	z�n7z#�r+2��Ҧ�w��ȣ�߉<$��b#rw�ӣ��։�'�m�`���,W`��ɔ��r�X�͒�5'�	�X}��(m�Y�&�v�����1EG2+ts�yl[�!�;8��0V%��f�Vs�9J��j[�������@���巇��%}%�S�?���K9�(�g��5�	���|@���:�J�B/	2�%G�1[�k3+�!��4G���=�@F����Rᭁ�Ա���!�ѯ1�n}�`���*��]n�Ku�;;{��FA&���.P��S�I�7��I������ഛ�4J��w��H��j��]�����>DY�f���~	|X�%�C]��I�2x���|x�o�iI���ʘ6�i��Y��j����m�W8�޳�rS=���Gƅ�ݵn �����3g�7���Y�q����,�Ї� %��7o�J�cVQ�7���ލ�U�{ӄt�Ǐ�'�4y�WKp�-�6������ϴ�H��Tlw�C2�I�Ǖ?�]1a�}�{���L���_��a�plZol���5�޹�pQ�'�`����`�(�9p�A��}���N7�c5%��$��a"x1�Z�q�_��3`F���f�,ow��y1|c}�1�/%�n�\������3Iz�4�ρ�c>�с&S'�s�������m�qg��{�N�P���l�|�۔��tc�?.a4c ����z	�"5��B���G��i�H��LzC+���d���=��$�&�����q2g�j�ju��u6/�������J��f�"x�(�L/�03�S���6'�4�A n�^��̳��o�fᠶ�d�\&�G�9+��m��$>O�O�/Е����c���Y��T�b���@ܨ�f���T�t�xl5�s���g����#��'B����ާa���ȧ�]|����jQ���{{��ad�⤒�_/���I����ϴᙻ�}N۔D��j�{U�T���-���B��U�u������ ��@l��Bm�
N�tVX�1�eCb^8�L��}�2V����ՠ���@7U�L��\s���n�&a�n�����FX�\7<~�1�kZ�;p9A�)��k�1�33��`�|4
pX�IC���ދ���<].�	��\k����Z��>�����A�r�"�`N2�7��e ���V���O�ߊ�T�(:/E��C��sd)���Tb)����L��o����wi������qI���M����}�T2��S,�k��"ߌ4	�Y��/���՝����V�$�&/PRS����wuQ<~Aŉ�/]5��ť�oS��[;p\�w.[¢؂���W�L@6���T:9��mRLKs%��v�L��vb�8�q��K Ԑ�����C�t@���<<�8֨�ՈYG��ȹO4��x���E���]H��^�e��[��1����!P�9�Z�U]�ho�&*��_��7&������/�w��%�{����ц�g+�cd�	�+@��ܴOȅ� 勼��O��H��,yT��A$�ߜ:�f����4�{}	#	 Ax�?,�|D��lm�?�.�\P���J�V�s,��	��}	i}3*��0��ĳ��T`�Ʌ�+��X��l�ѥڐ�~��c��v��W
�fЉL�]�m!3�{z�R�Ҟ�M��LE�KWَh��T$ �c����p`ǊR�������ĸ��.i'���t�g��+t��r�<�rj�t� ���q�ל�2tB�0��D�SwKa�jе-jc�)�����\WY�܂�d� ���I�_�(�	q�FT�>	�Y��]3����.�WxWW#���Y/���2�)e9��<	��̀��t�iĬ��2Ryu�~����g��~��:Tf���b5�W��g�OV�(46�,q:�T,XO�(��}&�75˱�h�ޙ�7�'�0F����������n�oaho�DwRjd�(B���{`�;����k���f�ެD;isB�һ�΂�N����E�8s�� �Am6�f�oE���T*ֳMݫh-KG���:.�|��V;����-V���1�]t�)��	*U�A�O�||6��?�'�CЀ����X0/5F>��~?C�:q'P��(9F�v2�X�>#U$��� c�ta�8���"��d(|������37-���9rb%cF/�V�J���u��_�xk�(�"�wi�4��ֱ��>}�>��4y���P�f�P����i���`�sS�_Lމ�(����XHv���)��ڕ��_�����3u����J��(%��ba��i1q�<�%?מ��kf v�t��_{����!�ֿ�袯�Ԕ+�,�U�Ul���"�\)��%���T�J��^��%�t��E��͍����(��9~������"a$x���![�ƞ+��ȅ��N�Rmv��c���CV�-R����ӂ�Űe�,�R��t\�3�m�|��0Rn?�l �x!��Q�;���:�T�f1�	��3�B�1�<�J��FZL9�.`'��H�Û��Ovg�w��}�ϱ��s�k���h
g�?�G�Wə�
|ˊc�w�p�Ql@lG��e������v�0�Hx��C�'�+��r�R��?2ù���͝�G4my�鄱�'��n��J�M��3$��QfI4if�M�� ~R�2���'�7m�ȿ�^��������4�.��ٙ�A�GM#"�Dk�����҄+l�hZfG�L	r1�&"u��3����W���8��"Vm�~S��DM�w��[��Td;�o&��41�7+�iﶍ\?ǂ�2����@-���D.�u�Ϊ%.�n�AL� �1;��j��'ힴ5� �u���x@�N�w&;M���]QJOf�}�<,��?C'��N��cK�.�ͫ�*��00�q�Yxy��d���b��k�ƿ{��p+�h<���4���l�����!�f{�7Gǀ5G-z�~��8�	�^�rI�L�Ku�H�	�ӏ�L�̏Wm�4$A�3h����@, c���;k��k �ʊӳ�ĳJPT;��k�z�[*'��L���Vċ�K+�v�d�1���<��6֯uYTf/o��ܘ]_�9Z��7�$\5�5�a�=c��� ���J1��Ot�k�6����"�Ot�ִ]�u*���5��S_-��p��C5m�D{3�u�ɸ6��Az%�u�̖�f4�_|=����(�/tM'�{�x�	�����t� qL����a�4��9�5�!w�z���F����9UD��@gbx��\�.^$G�'��/Ĳ͋��H�"��P�d�2uhiS&�����/���@O��%�4���O/��/R�:Z�B$MS9���v]���%�^����������d
�{e�,[U4arc؝�)��Ǯ	h#��H���
�����I_&��Uh�Kh���qM�S��60�Z׆�ʑ��גR�MV��Ƞ�!�aF�����<�����M���m(c���~#���Ǵ^��5ۤ�h/ݏ){w򵌫������V�,� �X>1�,FP?���p�9b�i�L�yeī6:�3~�	�Sg�7ǚ�ËFY��[���%�x�>���c��П�m5�j��՚>j$:Z�Эs����U�61Fe��xfdh�\� �옘����zdvtg���@C~�(�,�7\�% K�#T.�~o�� �l1�l.�#Oc�`�|k����yM��)	e@ѳ��%��#�ڧr� ��h�9(�g�����v���dAQ�� ��adD6(eS�%�`Eu�;��mF��];�:�ȕ)W�k�� ��S�/+6�p��8�	��,�6�кE?�R���v��+�W%�MNƺ��Z���^�=���p�lhY�N�!���~tB�N�UnPTW����C���/	�i���/�a���+�{�Tm�����r��C��w@Ȝ��Ҙ��-j��5ų�w� h�=G[J��"{68-�x)��/���s2��A�=��^�0����h�'v�nn-�����0Җ�6Zv���Է�2�)���%�Q��Tb�0/}��^u '�Y$����V�@Y��������:R�}�M9���X��܈����O�nM�=�����>�p�b�|*�-�ޅ�z��DH��N�vc2�W9��=�`iGK�y/Λ�u�р��{��z�? ~	��Ac�~eE��*���7�UΤ�մ1�h5e�	�3X�C]y�^6�u2���0M�F���G��uř�=1�S���'�S���rA���7Ïb��*;��9]��.�1r׃T�i����8��&���15�n��T�1����%%�Ȅ���[%fq�e#J_!�U1��m�+����XZŔ����ƉD�����A��<��9����-9|�����]�cR��N�)ݴ�D�P��$~��W�[���\�O�􁹉���UFr7j�z�,:.L��������[�����HTJ�X�ů�\Oۏ��$'�QWr���Ç�vx��MC<��>���)��D��f��0u{TC��.88u�y]�Q��5(;"cHHv�IFV�)>�[�t������;p�0�*�i 겟0� %$��/�h(�l魝ъ���F��+)����>q��h���Z��s�����ei�;!�*�49V��������B���N7]=@����x��9^4�Y.L߰*��4�R<��rS�)X�o5�I��k�8"�p��5��Yt>�Rc7���&��e]��-<��{P�m������yqa�4$g�Ow�3рˈU�n��s����o��v9��53P�V�r��n���Q+N��/�f&�7�,7����}�ai;�i���wu?S챺���׳?H��[.�;��}���ZH �LV|~���X����l*^�nj#)�Ə�y.�N�*�%���D\ �Ύ�cSe�{� �p�S��x&�֪��{�Z����:�m�^����N�?K�}�Lv��m�\%Zٵ�i;x�j��jҙ8��D�	��թ�r"��(X�7����Kݨ�],�\<>܃���B ���jB6� ��>~����m��֥��:�-OLf+Dل
�<��
P ��G��R�s���6���"�J\�g�3EgZ5���ۻ�Y�@e�b��)��<q�'X�GHa� �졮�p�ݟ�N��3���Y�� h�թ@�1^ʎ���g �Aw��^��{�L�υ�.Q�w�\Fa}; ��&��&���2`��9�F�$��;EY�#�Ťc�.�'�z�J�\i���1���ѿ�?Jن�F6n�d\(4����y�����/%?�m�LT/��n	272NgQb���#��~)j�޼����r��P��Gk�`�9�,�r��(�~�ŵ�Dt}��3��Œ�\��)G=��F�MV^�~�r�^�.��� m�Ҟg|6[�@�PѣQ�M�]-/a�^�tU���d��uS�;n�t�hC�y�S�=�]�N����y��ߎ�����j�k�7ك#� �̿+��U�*-�t����L��ۆZ.H����Z$�}�lPe>��B5ZC�:��`&��0��P�50=�g�6��S$f�i�	¸J�+���:�f�z��15a`�Pʐ��0Fh��6Åì�d�~�|�6���K���sR���CCZojn�)��"(�<"��NT��	0ջ�
�%[96�(ʞ3�T�S���;\�jkqcU��R[پ�u�5r���Tyt�D$5�;"�i6r{����NU�Ӹ!�C�]�2 �yx����љ���/����XLWB�r���K@Oa��<sn�ߢ4(KW� ���Y���Q��A�P�C�-�H1�����U���M�K^��#g|�y���9�7�����E{.K�$�@ɻ��]3{C���hS�<�����M�]V��5�狏X�� �v�h]7sC����ؗ!�Y�������14͍�H�P"o��)W��*�c�#M��u�{_^;���םn���ǁP~2;���)�.������z0�PUC�{�5\��hV�m�~!/�즬�N��P��R-��V>�C4E�~�YW�g³��kۍ��x�~��90�G/eix���S]?ض����'���q?{TA��yCE]�Q���.�"�M5��-U�/��l@�m_p�B�@	�]�d�>��6��k#|SGVyUL��I�����Xb�_����v� �-��q�.渿�h$=U"��L�唰Ҹ��Ɛю�p�׆�͊���jm
��Qq)�u�{R�O�R;'OX����J	~��A	R�h�0Ճ�5'��Im�A��bZUfU!��{�/)�{.��r��R]��+�H?����	wt@��XA��g&�r�.9�=GԒ��bS%n|g[| �J�wX��
V�Ц�3�)�o��? ���D㧼;2��!<�p���^�_�RU�ʜ��X+��)}��daG���	���k��3�ͣm({F߉B��*���H�߷����W��m���v����E'��r;[���xg��H�`;ɱM���&NB��ȓZ �$N��F%�?	(4��e 
G92�:b�(C7je��.��P'�P����|�䋁1Ǫ~�M�H��R�V��' ���{�l�C�pi2�X]���=ѱ �u���ւկh����S��1��ܑ�v~�]�9��9SO܃"��u�vM�Kc��uO�zk�k�e�i���uye��NǮy=�p��F���4�l=�ՙ���Spn���UچɅ]N*Z���9��13�V��'Kt���R�,pD�����2j��N�L�D6-�H�"(�����;�-+�*� ��`2ѓ�E �����@���*����^[��=?Y���Z�'e�*s@˚�:YR�(�����n�p��A�`�ҭD��t�R������s��V�钐��x��r���?���|G6øÝb��!�b.������8�,Me{A��h \a{���_����	�VA-���gX����6�j��~���S}09>�?���8=o��eԾj�\ޫ9���Y�6�J���;�r�*ϿZnbu�	5i=Q ��%&B~䒖jp5��������]��oR���N��0�)`��r㊃�&;>D#��^F��b��
`K0�t���)%��180�Ä��ʃ�c�cܒK�D<T�S���ƈ��Ξ#N|b���@�b�&pɋ�&�t���@TFŏ�.m[H�.r� t��]�-���(\'á�2E�� �!!=�!H 7�d��(� ��Q�Ol ����c9St�m�f*��-��zJ��W��+�!w>��|�d^B�����SnvN�N���r���7�d�5�u%�[ׇ�}adoFݫ�4���P�����i�֕���'���r%�ݏ;O�P�׳��G�/�Q���!.u7��"XU�i�lv�_��\����ó3���*��B�$�A��=:z4��a:�S��N�4bl<0\֢l+�@�l�[�t���Nl#�Ip.DG�11rp���]���v�ɮ��Y܌�˕�U2);��jM3�[/C�E�#]�(�R���Ym[�v����*_F����چ"�c^��F�T�$�YH�K}����y�H��3�Uu�*1��^�Xj?4p��'��w��|��h��j����[���)����@s��n����=
�O�C_hsj�@���M!t��m��3ŭ��xpk<��<"h����\��@���u:�8�v]nkY�-�]��7F:���LCZ+�`�<�H� �ռ��'��X�sC��͇��{5@�n�7�2�u���n��� �sm���]�ȣϾP7~�=u}�@�w���U�� C6��"��ie�t_� ��gx�-��v���f�x.�a����￉�+��5�?B��C2�)geUU�S���*'�v��_�tEȯ��d �����4c�188�5D�_����>ŝ�?��JP��pj��X*���H��22���µx��mQ<�{ϋ�w�V���tUݚ��վ�;��m� ]�;B=qQ@�`�xr��pA�aEn��W�^Eh�����W�=k�^a|K��;T%ˑ�z}Z�)��d/I���u\;�~���ڛ���JEc��ADJ��R̋z��X���(S?�@�Y�J��Ґ��f7?ԩ�	��b�\�Q%������8u�'W_��ظS��/t��X/�2��#O�V�8T�7�H�4���:8�.�,]/�v�`��S�вI�J�s����ot-�\ڤ����?Z�O�D�#�7��d7%q�O����x�`��lV�@(ދ+w��)����}A������翸�Ҏr�V��*�H�֪���1�0J۴wzt��l}D8Og�����7�A5�.sC��Fiص�8��j"[a���^d�%��r9s����4+�Ǌ�D��mhv*��x�y<����S%bAL�3��)�N�����H
Ag�^&�Q�O��_��|�g=���h�t����m��`��*�A��o�)P��1����7�ܨeh�;���2��V�J�A�'�EwFP�����^�"��op�U�izH�Ii�׏���.l/��K��K��H�i�N�H��I,���}��c/z�a�����gB)�V��
$��9�����jhT���0��˷�5�X�,x�LdW���L~�+�9�z�	�YP/d�[�R+�|)E_���Օ-�z�71��
�2�80"}�	%^�H���6O�#Ue�^�g��M)��B�c�b?����|b�?�,;X+p����~̍����K}�)�[���)��������#_���!����I��ۅQ�ۇ�A5�̨y%|(2y)Ik}k{�=�uF���%L�H=�b$��(i`�N^%ǮdQ�JA2`�q�+Z��$��^>T��I�
�mj�U6��b�/E�o��؂�[U*@�+p�Y�!Z��?0�e�w���re�Ą�k��wN�E
6C��&
����@��5l뙂l
aR�rn&K1a����eɷ���*^�w����暒�~u<�ˈ�}��^�0�eO]�i��#���0�VF"0��7�^�/��J~�<Lh�/3t�@nZ�%T��l�� �!�o|�t6�h�K%D�}OΛI[���'H�ʚ��h�U��Ӫ��-�lD���fy|��䤮V�s��	����8n*�g�D:�g�5�97^���^K �v�_kGj��
	�l]=#ST���'��VW�ϣ[���V6#��������Y��=�N��d��^�}�|F���{�Л��tg�K���kc��ʻ�5��5�mŨ��|���79�p�G~Jx䳴?��}�i�-�w)�ǔ�lL6��x��Xň��Bt�)(ɶh)@dLx�=��u�u�vQ�FdS.�Q�=�0��1&d=(:af����}*٩x-�i�-��f�	�??=�왪��U@.��V��b]_\�&0[�z�L�*�ٗ�ĳs�m���T*<�NfV�̟%�Һ*-	V�f�:���?��iB&�r-X?�=5��芤BO9�Un�&3��}J��Of�6�>m�[�2�&��ɹvT?�2h�,�2C�!3�+]yȄ�e;��� 0z���}0��&E��#K%��gS�N��L�C��8pG>�ÀD������]�/^�)/���C�J`z�kw�g����I��6�7�I��*Q�� 蹽��q��8���fϸ��j-\�u1#��CۢƔW�a�m"��>h�j�������l*7�ۛ~g"�4q�\]���(��t5�2�G�~9:矾��X�1�olT���^� J�;H�9��J7Q�m�.dhg��u ֱ�����ba�X�3 :��	iOw�q��#^��pc������q��׷��{��s�)&�$�|g^)�֡��O[�XAI�B �rh��Vvl��ڎ����5K�_(+�r�W�=����<ٝ!e��4Wi0��� ��P#4���]X	��7W�u�*򜒡����� ڨYk��|Yƽfff%F���G�)�Œl`,�0�;{ ]Q�5R*=؆��t��)�W�$�$0~��ʡ���P��K(��T��˲K�>5t���U��t���|v.G��z�L.!,�GWt֖��J�i�Z��<��1A�YF�Qs~��E�˄5�rB�>o���AXx�������Ÿ�E�r��5؝GG��q�V<F[@���k���>�2�5e����d�oj!$�2�:��x!�rTq7D��E�E-�߂4�<��G>ߩf�S�7S��^���Τ9�ƍ�x�7���BI��tXV�l�ϋg��D�ͻj���}���-ʒ�kޒ��{y#���SS�s�W5��]S(�������F�|/�ׄ~2��˷4�p��i�H�.V^wf��}�p~2B8e�ƚ�{�m �
F��Y�WeuT!��D;��-}��m����L��J/�y*S�ዮ0�I�,����C�Nh�H��\���fOئ�B��B��4��~-m+�f��4�r�i�|*^3;$��M@��e=������jZa�׌X6���3#��W��̭�g(4��}j�<wrK��
�i���^�WhM$�=�ʑ�,��'������;�w�J#^�o�>cq�k�c���|6�#]�-�EJ�S��x^v�ɹ� ��"��8��k��e�E��3C��������*_�2�Nz��!z���O9�mLY�K6�� �C��4#�H4|wtě�$m�ܹ�O��t�=��H�V�}`e�����E�c��he���%�J���Ԑ��K��or"9O^�
G�q(�^��m5��A@���a�:R�,�i�Ӑm(�GbtYI�M;��l$��%��I5ˇ��z�����4� ���"jYuMd�jƲ��[$�B����G����>����8t�CvkA�	F�Ϫ1݆H/tl]l���1l�����{D�#�����5��9�;�B�z�`ӗ��Ƣ�$Cw�`,��a�]-%����0�7s�Y�z���?s�}^�Z����Y�/�R�&Z5p<OI�L�T��%8濽Oy^@���5D]�F��P�;g�G�Mt�@d50�����[*��S��q��`�n��}�Qy;,r`��@#�_��R9r�z)$r�"����nZ|of�,Ne�^Մ)��j�uW��*j����Y�8���;��/�M�1�g�@D���6�:!�<��Ƿh�$r�'��w5ŕ�o�a�����z+ �v����Bw�B���n`C!s��n|�˕�(�ЫO�$@��x|~d!���n=ԟF㢼 ���t�gנ�hez���_ �	\%����P�3�P�˗B8�`���}�EBr(�����Py�&yT�8�`��j)�ݒ��7�R��\=���{�H�	�s'm��Ƌ)��o�u��)�U��;2��䕱���Btd����Ci���Zē5B�#/k�߫��=�gv�X��S���wW�Ark��<*JF;�P�l Ri�	��^������/a-��S@��P�}�$�3��?D��ޗ)���^eU��k�t��F(B@�ƀA
��n�I�m*�=��k:nDbo͓g$�FU�.̲7@:3��gw�Kq����N��a�hx��,��\�P2��p+����biu����#��*�C�:i�T���#2������OEl�Bd:W�_nt/�ET5v�
���bxs2�䈩';�i�"
(���f�}m5,���@J��V
�q�5�5@9u������o7�Elnh�6/��S�0����=-����D"B����"E7�����D\��Ī�lb�^��KyA.���i���p��������!�856�	 W4 ��� ��퍧�d�i���m�s�Ј�p�i' �_Ty*�� ����d�s��������b���a�IX�n��i�t�P�F������a��A���)�-GV�A�L�txj��\�|"Zͼ�$���F{��<9f���5�L��k�̃���Z$���{�T��_7E�*<X(_���һ��"�O��F�̮��H�r��2;���6�N���Y�.�ո�|��Ú>��T�`���~c,+:�T�5��uz��3,�������|}�l�IG c�K���SV�H�joyC �V��R�$MZ�)Ӣ�U����'��6+��!#�)W#Z��SE	1:����iÂ2N(�:y@௥1$�q̛��yej���J��ehk4�=绵>K��3*��F��s����w�	*>X�b�D`"Ւ$o4�-ⓓΉs��gC��}S�W�4J�$L�r̦z��`�'�tY=�K]������b����`� z,�/T��惞�Qy����i��%����c9&%JQ�R�K�2�@@ɥ�{���[�`I%�4�?��#AS�$H��)Y������l��)xt�7�yU4�[/�[+T��n*� =ؑ�,������G,�R���O�4/��,Q��E�eBz^�}�*�,"�ٸ�z��S�z,�z-�������]ǐ#����~Z �4O�-SH%	��kI�Ϧ�8گˢ�0�)�ޜ�f��Zͣ���� �t"��'y�f�1��	�,����wǇ44I�����l��3�W��|A߬}f���ǿ1�q�ȃQȖfq���F�@ZXx�A��}�@�+��wu�C�*�?�Ee�ه��h�
b��1T�¬�.�������P`�?q�L@$�-I�)���[i�J5�&��Α��m�]�c���=�o�_�o��%s4qp�Rq���2G�K�)g+"^�_z��E��0lp} �4W����c��D�v� ݲ�Q܉���&!��se% ��F#`���deh�]�.�����ha���O�O�J!�-�܍)a�2$��,����Ì�9��M�g�ą[0[UTK7��h�ם.����UU�`΅O�Xn�YI|�Ɓ���o�8�&��;:�k��q �� ���,�Ǫ��.�c�Ē����'̅����2}-'�87���s3�%�����e���tG g�ɏ�iE�9}C�U¥��܃sK�lN1�Qp&�:��Ѕ��`|aٚ���b��js�7�#B�i�H�bM]d�x>A�&_qWB�����f��~K(&�\����nH��(�bX��w�`�Z�~��M�㡖�W���D� �b�L�&Q�&�߻A��W�[J���8tB��s��	S�{�1%T��茌	����ۉR*7��p�3��ӝ�n=I(Ԟ����
����/����)�=�{G�D<<��=y��7�;����m��Qa�^�>�n7Fح/���\�' ���|�� �(���6�wu��5��^[�x��_@��n��I�G������h�r9�_ jW�Y�����u"�7A@l�a�pUϣ;�5v������zv���?�Ear�����*��#�po6E�"뜧{ڳ��s�C�dz\@@!8=�H����oR�|��e�u�%��2���Ŝ�o0��������F
�L��RV�_�I:��y2ݳ��L	�L3ذ]F�i։tɢ5.��u�4���-S�5��-]!�@~��k󑋘3tS�!���?HlWӘ;�w��1\ȓ�����P"�M2#�j�f$�1���u]D��t���X���<qjD�JΪ�*D�eS���h���۞1����~6VG y��	[ *��fW`�T��o
�4FO���M�E�	Q;4��ٶv>��|�����3��0c�t��i��ƉR5��M���v�t�X�W$�g���|�&ƙ:	r�{r��q�fU익h��gҙC�$-E*G�BL�H�S�⭔�\���V��^�}�'H~��"��Z�u����>[����G~/�n�ш����b�=���F!�>�[��H���{˧�I���@�0a��y_~ZN�-�X��h�gpj�X�By-lC�t��U���s��Ǣ�g���/0&���axυM�\h)t��Z�Q!>�L�2���u��y �^�j�3��5��eMg5N巐�w��֩VK9��+��\��.�ݐ|S�Uz�N���W�m�,!���sn�l��t�e�8�nw5���ߒ��F���LPy�4K���\���jm�ᆟ�����b��S���X%���s�Cʯ3�~�x��o��'/��h{�c�Jτ�A�$d�P]83�\S�o��V��V��kg�$3����f�ẻ����sm#��eOl
D�H�U��I~s�>�JQ�Mfv�0�8@��(���	�i�0������ܷ7"���rֈ���۵i��5	����~�w����Edm��|YE��+��=��=W҂�K��.˳�$|��Y�Wv�c�	^�U�e:HR�li��F;�
Z#�����S��0I�Y����3�t@2v+$�sE�i?<��]���Gaa1b�!���E������.�O~��s�%2$=� Vׄ%&��"�㻤FD��/wW����3C$�ٗ�-��d�3�2�� �&[Q�z���4�50���{�A��&��o��?��=�Y�M�v�$iE\)܅+Y�.z� D��߄�*�I�M��k��$��Ԝ(_\��WÔT�#F����B����� ����Y���� o�CtskN�q���&d/��?[�|ch�n-�
����@��>p],��.*5Y�j�[���h���Jw�}�Li�okR4�\�[kY8�P�^	>�D/m��6��Ik/ސɮ�<��[$	`�B�����q���eM�m�y��i���}�6��Dc��u�� L���f��X�{�X�3�ςw����K"JRa`7���2;�p��%%���%���4J�c��g<�l��5�!ZA,>�G�Un�xù"[�Rs5�."�U��QِAW_�}�Fe,����	5G�H��h4W�e�{���7O;2� ���h��T��IѺ�R���2B��M��T����|x�3> �DC�� ��Y�c��4����&܀��?���*�CQ��8!]�771B����Sqbw�c�[Rw�v1��TCX4�����l(O�N�=��M�2t�}g�E� zI��?�9>*�����-h����)[s�w�ѶiX�pu�M� �*}K[[Dfr��v�1	'�)��1З4E��;���P���P^i��P^�1�>(d�HJ�&7zDV��s�7q_iW�I��x��=�$���i��O+3A1(� U\�t����R��'��-�'.�v>�T���'�6a��Vm�Ν��j>�_w�ME�HȈ��*�؞Q�������ص{%�i�v<U��ln f~$�sa�9�<_���[.��aU�S�!�G�w��7�o������XR)f��h0aZ�@���ɨ6{��G�|c���y^*1�U!����[_l*���ZS
��yl��Z��0�-�њ���	�a��be`X�����8����)4��hq�ɍ��0ƭ���q�:�b�X=��c
��
~>r`v������Cø�&�v+��E�Qk�=t��E���=@׸��T��0��Bբ��;/�(KG�?}؋֦�^
6g�-��k_lj�uj�ȍ����|�r��r��s]����ԎeH0����;Ƣ��Z��f_��3Et�2;�O���ڏ̇H�W����NF_�-��_
^$M<�g֙NC��������F�4)V#E~��fֆ�|W�+�Q%�C�r���T�6�4] ��"wK�B�:�CH�#Lq?�ٲ���
cu�E[�mo�1,﷌C�EZ�}L����N!�3��~BJ�[��s���Ͻ��B�6	6:"��'H"cq�2L��i!A�o�e�fN2�3�����u%��|$	v���B�ΘzG�I�%:�30�"�R%� fࣿ�,Vz�\�V��� :��r�p��	堄ܖ(��Q<wQ�hI�)��[þh�s<�����&.Ž,$�.^-�Lԑ"h�$�@q"H�n�U�_=�'���b�T��B�@ԡ����we���b��tA+����v�TL��T�'�ަ͡9��̈́�Av=y�����pg���A�e�]c�dR��� F �1Dwћ{S��20�`���K��n��*�to�-Ds�_��ܴ�R�sѡ�?@�G�.�%��Dc�n�r`�z�S̷�8Z=*�`���\��ﺰ�����G��ة��cgp�it>j�����aH!����@���@��Ne�N���!���-�?�����%�,$:z̳�~��u
�=�x��U��N���+$@�y��X���t��w@���4�t�E�D�j�@����Kd"=!�x�mv����S`�d`J9�����N=���%y���:�܉�J�_o�@P?�2�}���n��X�e�)�8p�%��S;�?l�Q�v�,y�������륎�͞C�"ث	�U�uMy{B!�p��W�%?�c��B��%�U�>eV)P�~jMpq���v��o���X��5�#@��3S�����<6֠6�H�o8��SW����r��~υ g�T���K��_x�$��A �I5eO)}%�}.A\.|l�e²�gmqU��8_�ϋ$4-��$W`}�/b�A�l��'��G-�&�j
��g��s�U�1�����|򁑽�./Z^�m/�2�,�?��Z�`Z�^�7�6P�Gg|��}�d��K�(�ܟ�6�����S���U9����s�tτ�Ե2��>v��̏����(�׼�0��鍱"Mj�i��+猺����
��.y�<�7���ۏ=�ASDR;@h��.-���=p�Z}
v��M�F��$��"��E�C���l��!�n�H����<��F+t�_�Ty��ά���{ X��w�x�E��+����a[��iҕ���s��u�S���+�Ĭ�071���jUB�� _��9#n�8��7�H��y����Y��(�_�*�,pe)�5'Ǉ؉ِ+�8��4PI�W���s�ݾ�RQB�t �B��9�[Mg��������y���f6d5��M:u|e�+j@ɮ|[X�-��J\��`3�I��c�\�����M�����h[ߩڣ*�1$�k�!��e
�>��Qw�e$o
sm��'�Xh0۴�}G?�py�R'�����]�2�ӭT�1��e�y�dQ�?{�lւTG�Tj�i��n�xϪ���B=M�԰%nQY�!bbc��wĄX6�Xov�`��A��&���>�;��8�p�5OJ,��L��j�1��.�X+�֠,�P���t>�Z�t!�?��ĭCi�|S�2A�Ƹ�Q�!�&v@xX6j�0�^!A- K�
-epR� p�&��׽nH��EH��������A~+
�[W'�j��fA	SikXC��M(���hr�4�/��_��?�J�W�,�r���!;�SBiN�E1l9r�kK`>�� ��2-�K�~	y�Mٮ��E����#~W`�, s�Ӂ�F�"����$��n������\ �����i���p��K���/� ���Lg�~�P�����ӬR�j�4��S��L&{�2��q�D)�x���Q���gĈ�����[&@�����Po�����ɋܒU\Q�\!\ �r���+��~����%y����#�F]��B�ݥ{5�;e�)XY���?�"�u)K&�!�����#`�������sņu�0vRH�r�����`ۇ�]�*bԽhŉ���^R<VoFŨ,Z�u�G�=��h�We��K����맓R�zE:w �>�&�=��M�6aͦ��i��C���R����_�Ӻ�'*���	﷖�t����ȃ����Hw�߸��/t�#��`]�� ��v\��δ�􎏋l��6VΌ��4x6�us� ���q�F4*��Tj׵�YWjJ�k{C~��:�)�H*)	�z-���)ԗ9�>��?Ϛ揽�4gI�f�����x�s�k�BQ�75I��N����S�Ms��OQ���(�"E��XG�S�W�NsA[Y���I(S�<B�:�6	U3<���7"T�n���k;�9�X#G+�C��6͛O���u��N^t�Lҵ?Q����Ƨ� �ؕ}��#�^��l��G�Ȟ��ϐ�7-��U��J#&�t���C*�_̹��s�H�<�����g�v�:AL9'
�A]�7����1��	�h�-�v+K�y����ʏ���G,���b�w?�Y�W���������P��n����ԽK��&�9�BĤ?�)�)�*C�?�����V�Tꏔ5:��a�'ג��*��s��u+>�]��g�nXޟbs�`x9Q���ɗ�H�Sm�g�G�A��l��X��e.Mŧo)���'�_��[>S넆�;����W�>�c��W�:��0�r�OL�ʠq�r�+ۈ9�
�����l�����?�k�#F�u�Ճ��G�O>���Hl̏<�����((�����Mf��<���3����<�{�!a�+Y�iV���Ǚ")D����/7��������m�LΗ��/�_�n+�a�*Y7/\_����F��G���9b�})����8��� �V�}�/ë(:�	�4B��d�p�4n	=� �Ͽ^n�������f�M/WA�*Ы��m$0.K�&R�tG���|A�� ��%�-�Ą�T�u���C���K�)���%�M2��;/a�f;.3Ϧ�X"�n�����ƎQR]�o�1����Ը 8�� �{�S;��e�oѦl�h�+�����F��) �=�k�P���V��v-�5ԩ�
���@�Ʊ@,89!��������6�.��-���E y<S�⚠��;�L
�N1M��V�C@��m{�~"�˜^D����'�U�}��]�{�;g��"rk�;��Z��t�`��ս�u)�<����4|�9�4��e�'�u����ɍN�@�V"~"�sGz�a�ؤ�����)��H̪���|.�3^��f|x����D���gˌ�
}��@�� h]��T�h��@���f�g��r��5��(��Zqp�R�ӹԵ��J���m�P@Bԍ�Al5*����2�Ǳ}~!�a@����w�(<Ӓ�@Q�����D���!	����4ʎ�L��Ea��8n}���8����}2��e,�PV߅н?�s�y[�Ya��?���z��p�iQ>�(�ގ4P>��Z�	 �9q�:�t�:�Z�x%(���$�
�R�=yZ?/��h	��Mۅ4�����U��ъ����q��a��mS6B�]���g-K1EQ9TWU �b��n�7s{3kԥ)VN��q�T���*As����6?��w�����)�������QK���`�i� _y2�,����7���qmuz'j	;_���T�cLK_�,=S����t~�!LU�9 �wq�\S!�e�[B: ͅ�v@E�������\�Ƣ����H�3WB�� ��Q��u,�7�6���[��='�0��A;��t��nm��;U�^DNV� [�o�e�(��"��9���
�L|=Ji��Y�M�T�Q�|T���dr�TD�AU/��Ru�\���#�f}���v֞�mL8;��rA�/KR;�y�z!Ш�c��^��0�_7t�Yi�G��@ ��[AVc&��P�r �ΰ�?�q��#T��6GrFu$���l�^���֩�9�x�G����5zـ���|&�M�Yp��r۸�BF��`g?U�����U�[�G���Ɋ
N`z=��\���5�>�vV�{PG͉j�ՌR�0^f������Z�@`}�h9�����D	�ޫ6y���,o�}8~��0��/Gx?��l��"��K�����M�:(� �s��M+�	t(s3�bn&��Ȗ=�������5����K�tYLj&�Ôs]
�A�;�Nw���c�F�σy�`�mX}=CyN���EP�á1n�:��񔂏ܳ���6-��'��l�"`[�ހ�a�4�`h�,�:h�H
Ȳ�f�$�O:,�cvK�9B��52b���O���=�����mw<�ʕQ!�"=d���9�0,�T�$�q�Su��ux6���_��G���=�DIP09�!B����؟��� �^��X���i�Hm˨="1g����\V͈�y:d>��uh�q@&њ2�U�B�D[h�N�M���0,�%}��C��,��9��GMό�Y5����!��yu�7�N�O����-?M�C��?UB�_�ɤv���E[f���Z[H�4l��:X��ڂ��Q��J��Q�� �;�'y�3�F+M�)Ey�ј�kq|Ĵ.v�KF���?��ܢ�e}y#��<���֎�]&�fY#><g<g��8�=��a�NH`�̾ݸ ڿ�w�9Z�%(p<���E���ХM�|��Y_���ɔ>+����"���KﵼV#J��'_9��#��^��O΄����T�O�y_��EC-~^ҫ�Fx�|��k�1$"ܶe5��*T��~���֙I��f��h$�x�E��)ǸIK8@�����8�$���V��*Ƒ�D���4z'i7�"�՝���3�;JO��n���q���I{�jݢDP���=Wk�e����LS^��L|Q�*��He7��
�QqX�+i��[E�wP+o1#~WI��NQ��Ź}���;�PMoh����Y-�f�VM���{Ed�Y�~;��i�[L���}^o�ź���t�G6흈�A��h&� ��:��s4'����(5�56���aS��<o��#�?c�8���%�3 ޳�`A
����B^�uH�r�^�<���Qbb�*#����������$��p/���`mU�߹�3��N��0`\t�@J�c������tw��G]u"�b���Z}�52w̿�T�P�mr���_G��a 
 ���g�[�=�1k�	��R1��D٬Uܿ����F.��	��T�]c|��[��Ԥ���6{a��y�+"�h�6V�'��xaGgf���W�~Mεi�92*$&��v:u�M��X��-��12��H�6E��(�+ �1���R�&��v�d�r��C$9ڈɝ����$���9�:�3�	����kG_xV�f���u"	�XO���SX��Aٶ=�+�������Sw��˦r�'k$~)<�ɅEk�x�ނܺ��`,���$�c�Z���������Ț4�68{Y"4,�i�݌�/8��iuX�aYe����E�ǿ'6O �錄#��6�|n{�߃�����L�����0���m�10S{7�<�"��d�!ՈP�O�n��i�J6�8�U"6񤑻]z�װ��3�b�K�@-��b��M
+"9��wJ�n����TÂ���z�(�0͂���p�O���H�,P�la:������;g�9]��/�r�U��u��@u{T�z����އW8�9ѕ/�jl$w�Y8��;��UȺ��%	�_=��g�$�[�gk��$��%
L�@a(4�_���CɑOg����b(�PN�˞��ٰs%���%[m�[ml����W�ͣ�h2Q���� ��9��[#Mw��g��)�� ��#�f�-�+mqWýM]���zJɅ�8�p0ސF:�A+:L�f�`/T��@O�T!4%$-�'���qkl�I�|�jc��ˈ��G�\T�_�#�D�?�0*��\h{'%�~"]�QR�X��C��nګ������N���j�nm��F���j�Fn�W@@4a�h�ޒ)\�т�4K�E���� o�µY�vJ5Ʀjb��AQ��<��  �_*EU,,U�,e�s4���y�_�'�~�2z�%<�u�CuSm�N���j'�\X�@8��F0�V����&��^�:�ʜ�-�@���Σi��s)�Sր���o��޻��"(��)�ץ�����1}�+]�į�����_�6�&�BO�������I����!8)���.�+�g[R@�ʧ`�J���R�V��꥘�e���!�i��~߇�SH<_��Q�L]�PG���>��n�����*4�Bc��^N˅�@D|坱���F�(g�B���5f�a��]GSr��xc>�,�:'�堻6߮�D��z�-��9
4��8} ��]�a	n!pC�3�N�Cu�P���?��Gץ��\0x?���v�\[� ���J���~y��f.���{��_K"��NĹH֭)\8��K:�[Dx1����3���y>챍�W=�C �ۓ3X>@L���Go.1�-�*e��-��V(�LM-m�"�,�Aگ&�s�=�-����k4U#��	G�.G�tK�����F�;x�C��r?q2�_e1^����R��@g�鿴s�˾_�F!�� A�ԯLl�,e3�\®�8���&K7
�4��&�
��~�6.;�s��� 	Ny�Ro_���J6�6��*Lh�M�`���eǖ����9u���]N�^���{%�#ĭ���_�0�g8��*�h��z΋<{Mr�U�����Ҝ)����d��Tm=�6�c��1�=���UOc�P�u�,\[r��(��g�w�m�>��y�,�;V�sΆD_fL��{��f��a�b]���oj�v�0�6�kšDwH���>Z��b��'����.L�_�^v�kR
�*Nߥ^��(�섮�LH.H��"��p�s�F�;8{5��9LO/,
�������xխY���aN�����JXސ��`XM���l27���<e�^
�Z_`���/3�0��@��U�0�
�F<X�.*�T��m��{1�ؗ0&���F8��D��S�K�����u��~a�#x�].z�,;�~�ɋ�w���6�>��K�%(;#�	��i��V�.����;�%�~��{OWݧ�ז���:c�8|�g�y�ʭC�J�'��0i����wZ� ��>�C��Y��ĵ!�G2w�?�'�6��4�(!^|Ƣ��2Rk�$A>��������B:`���r�觥u`���`M���R���͡)�����'��J���w�]��*��2
扴�y[�:&�@�᝷�ĐTO����L�&r�������{�4Y��0���Jj`�#��]���(��]�Qp�4���^n��ŏ�*}l��ȼs2�j@�1gϜ��
}.�X���>�Rè<qZ���>�)��&O�Gج��9�v������I��|�#�������AD	�n��JX�8$b��@N:[xf�f�2�6ٽ�چ!I��Ry5�_i0V�C���H%h���,o��nV\�D& Xn�ּ=��X	(e/]l+�׫,zo�؎�_x6k��N��n��٪}��>��,���rV�^�FO��kg�j��8��-�Z�x�D�;����F�ԛT�thrͽp��>�c�j+��}���g�Ӆ�P�Я�����;�(Π�Q�+c�G�%��+��xS<
V8X�?R�E����~��Knh�K��m� u����������^�&^P�F�\gp�Rqs	T֬�\?�A`�3��2�g:��Gn�~G��E}�@�O0V2Z�4@���E:�vo�?t�T�f.���
X������M�$�������N A�_���e�@܁í�Ct~ >�n���7��1���-�<W��w=u��]��#8�$����f˲�;� ���vSMY�
�I���"�U��S q�Щ�f�/ߌ�F8�zpĂߡ�=5����M�_,�DBރ9=���S�OmJ�T��ā޺Z���ME#\2����]�B�Y���[*$y6�I�t�� F�ԑĠk� �ޘ�(JWS�&0� �#+��{����'L�P!B!���J�#u�?���rN�8�]�^<�U-�ʟ��Kt8�pz� �����l��{�Q8��Ϗ3�v-�ظ˃����I���v�dF�� �	>��5�=��*d�HJ	�fC
:���aWN\i9�m{��
�d�zC�D�s�H��� +z���$su��$3P�$��ΫL�W� ��r��mR�#��;��̫9�W��(��m�=���� ��#��t[lne����M��6����M<)eΛY߷��S�D0u���lA���Qu��EY����{��,��Ǫׂ0���	����+�x���M�D)^�J����P>���ے� �5M#5�5Ϋ�<]�=ʾN
�G������MS�d�����|Љ��[�B�D��D[
��i�u�+-L�T"��ӥz ��c��e��v֥�Y�����7�9�7��}1�����4�L*�4F�=�UE��l	�I�I\H�y�`�O���Z�_&5ֽ�̹�t�A�X�'�h�q��-���w��0Okl����d���Xh� ����"c�Ϳ��?H�F	\�^Sxm���j&�H����%��}i.�%�my�(��k���g=K�ğs�a՜̵ s��F�y	�N!ު���d���/D7��O�����P���D ����N�0Ja�إ�ك^�˟HX����YL�퍛br��#d�]����o�}��v�T�΅�N��N�S`��"�Q�Ul�L١��q��!#�8L
�j��� 1����P��2��a+Is�\?4�F�|�*����֋�Ȍ�I͚�X���d��_����g��3���+��S)�jLe�K�4c�W���nh�٢��]"K��4\j>1BP����bi��wn��:͉�I�[�lw>��EL�yՖ�,'���w ��G��)|��5�����vg����B����� 	R,���:�\8���2(E*��/�G��b[�zM}��5Y�X���ȏ��M(�W�పb�>�4�.�fяH��c'z�6�]����C@��L�-Q���×s��.�� �Q� b'��/X��^Pz� $�7Ы	�	(���H;�kP��­���Kd�����泹vx�jX�s�"�bC���4pk���W����a����_.V���):�Ȇ�<i. �,�u΃з��P�<��QC���La�D�t�َ���2�W�}��Y}~-�=?�}�	�9S�t���]?n{i���F�t3+rU�v���#6�2�K!��"jw��8��+���!�|h�S���jȉ�c��:����&"_d�<I.���K�ħ&��;)ũ��ӌ(b?p[��e>��^���'vw��*gG�.�����D�9(�&�B@O�%�ms�l�����])$����>4�j�� ��� �H��N7X�Q5������ߔ4�r�QQD������l��F/*E�u.
�,]a�<,�9"�*�¬�Z�Yg�? �2�Ǐ9�9���	��$O���d�E�����;hݮ���S�<��F�E��Dc��N?v�ԡ��:��Ǹ9jg��fIo�]�
v�IO�F�w�A^2/�;ȍ"�|������Ѣf�A{�s���"�åP�4DX�Pv;��.N/�������f�!���t�
}*�������V>LW(FJ����%H%e÷��d�AzG}����7ҭ�T(	�ӷ�L����e pa��ȿ�b>�ȃ*#Fc�t� cH"Ux�{��.uI$܇���)m��;�,���-��p���y�ޝ>�?��BԂ��,Р�0��h��I���at9��bZ��d���/(,���ʿjƽ2�jXP-\�-Yi�i6���\���r�,Q��'�
�ܛ�{a̛R�>���6�l���m70�.'`Kr����(��+Ek����1@�o����%
v�εK;
�e�ӝu��Bqc��}0����vûx���&z1��k������l�¹�t��$bU
����]5�8��v���L�Q��$�Ho�R��Ĵ� �E��B����%j�1��J���w�U�`zȋYŻf?{X��=�U�U/T%Mt6+��$�ͶY	ꕐ�e,����팘,e���m�O!���4)e��ڶ�zPa���@?�q!j�M�	�����S&�H��
P6NN���u�Q�=ڏ����;�ܩI�PnB�o���q��G�Kj �|�����]�d�s<�~,r��+"IA*�RKD��������/
� I������g��%��n�j���Q��!*�X��(�ޡnC�ۧ��}_~�̻̐�2���g�v($b2O��=��oG��������[�驮2��@�Mʃ�:��0��AXC�JO�,!B�#�@Ye;$5�z���=�J��}��ذ#�/�	�������|ѳg��p6�l�k?���jV��?��j�10󸽒}��>Q�}G��#�N$�-�e�g\K�lB
�6�u$�Y��S-T�^��N��|Aٔ�X�U��B!9��;p�o�1/Ҧ|x�-����Dn=����|�Ie�OG#�n����ɯ��&��i�[)�4I�I�T�x�w�Ń+�m��Fl��_fX���_�V.k[K� 0�#�7��	^$� �����ܔ܇z�l�n�\+�Z~�)謶�!� ��z�������.��'��'�?�'(@U��}������#&X�/�]�+k�<����-w� Gl�
��ޱ+pSd;�{?:pTRF������.O�g\�&��t>)����Щ�����\9�!��3�'�(j���G�iP�N�6{�IT'�`���e0�bw��U��p��Y���5#�����3(���O$!*�*�Do���#F��D��^��[�4JW�h&9�1|�*e���-*&:���W��|���ּ��k�0*<ݪ�Ce��SiJ�
��j ur�3�� #E�WB4���P$Ӱ���(H�&�Wî!�>k��{�
��'���&䍮�;W�#W�L��$���0�����߈*c� �r���bq@�,���z5�O韫����V�H�X���΅È�N����Y��������9`O�=����Ѳ/هq�|��� �n���-`ٸ:����x���DH�(�*)�kT�D�ܿc�H7 մ�2%T��#1�(ϔx�Α�ֵ��:��DǵB�K��P,�?�HɉUl��늄h�zw��f��{��O�V�̟�/ރ��s^G|�>R��g��{f��{>:�wޜ��Z�A�<�-�]�#���q^��bo������Z�O���{~�ʨ��u�pU����>oe|��艈Q���:l��ok s��z*/56U��V�7�Ԟ[�W-�x��Wr�&��^4�P��ls�l�d ��O�aТLð�M}�f.I�b" ���g���8t&���)S����>AV��J�u����`d��c�j8(�] ���QC.Zc}�� ��q~�i��E%tL,�7j�M<z��+y>3݅�1��e>���e���+W��iP�?�8��!���pq�ak����z�N�����0ܗ�V-si��B?�V��J�õ�����ݯ�����~"�}?H�n79oR>���}�d�1#�������ς����q<��4�C�0�_3`��2P��e�j\�X�~��la���Ԁ�D�-M��o�Q��}��Wt 1��0"�U�ARͧ5���qץԯ�u��EY��}�&��:�*����-�<0�s	���D�����J]��3�ƛlK�!��p�� Tm�F?��7�5N�!f���@�9z6�!9Ewh9hx��HaR�h念���i��`�l~.{�Z���D��iOD<X���\�}�2�y����l�� N��˻���|i2~5���B�v빾/��@t���l�OG��І��z)6xW��$Pj;5�� ����<oJ�$	Z~"��,�I��a�����dU���8�' q?7���=\��Q���bu�xi�\B3~�YQ+V�>��^����u�	��Z JڬYO�k�c��|���e�0	�E�109����w��T�"���cO�N Y]�^�g$L;��p4ʢ?X�=�����i~p+,.��[����~�^r�Dxfs��^?����V�q�a}�c���	C�66�,�%��J"�45�(�v�<vu%�$����:����_i��p�M5��t������D�JA��G�{�ԕ/���ի������2���x����%y��$ڪ������1��OO�K��g�̷���rzH��@��]�,� �-
����Z0f��&j�ز�hTk�q���s{~_-��qf�l���������|�'��!E	������tRN�JC]�!Y^�w��%rي��1��Yp|�I���y��M/�`9�ڪ��N�����R��9�u�Tq�V�ͷ̯OǦ��0���o��H��=گ��D�٬�L�vs ���9��a%�ґ��x�;���$�P���v��^俫��y�L����jq� _:���+�A���Bی�5aP��5�������)�q�]��![2���oCp#H�/��#y��2�f���+ʠ�����
��y�/�2k��Y`�wD���ߣc�`�_y�o�b�Ҿ���S�LO�f$�G�t��ȌU߫ %�T��>p��� Csl����ޏ�]�y�ۅ��/h�ߩJԜ�������]����L�4� �vg'���	�
n2>m�T��oJ*!]1�{˳Ga��@o��d�J���Jf�p�/�� yY���Z�'� ��W�@�1W�Mc}��s�I3h����T�0��]��O>�5�d���V�m��j���-}������0��6ƀ�:��ל�̼�������?e��<ک ���-�T�L{<]���]b�������l`,ګIU[�e±�7`���4¬���2�*�A��nWt"n�h:�V�z�Œ�mD\ %Yp�����h�p�L/�YʊW�]J��ly�旫
�������%�i%:�wH�>p0�&��m��4n��&X!��)K��~&�3?�)7�]4|��2:k`F�{�P5Z`
�U&���~�C�uՆ����4�O�s&Ϲ�ÕR<���lBĻ�y�6�tU�^>:݆��d��hI.\|���� '�Mw�IK��M�h�˚D#O��F��Z�������Zd�����I���i��gS�g�(��� �g��^�]�G�6 (�P3piC�^ţgn����ջ;};��W��4����:����|{��|�A�Z+�5��bŗ%�EЎ�R�
X^�h����J7��m�<��;X#���$j9�r���Qxw�|:{�9�.�5+h��gR����i�eHǰ��:wI�����o�}����OqI��nVݐ��|�*J�Ɗ�NS �Wl	�`\�zɆ��a�a/�N�=Ə��0s�F����>�:&�*g�8��z��hn3�T8�Ow�t�«�����ɝ��O��@� WL?�Ӣ�X ��OUZv�����3�*��V< �r7:z��Cfb[�����B��1�ï¶�
��s y8��T�B�d`�%5�ة�D�b�
�g�
��o�;��֓��o�ٝ�1���)��ZU騴	�,����&Kg�*���J��Xn{IKe�M�B�z"c�[rEI庞�A�����.ީ�����` ���2ӜZu�!�U���/(��mFڧu�����{��y:jcjOd�W7����m�E��W|j��(�f���CP�N=�B�Us�bq�d�7]�b�F,i vy�����(f���d��XzI,��s�$X��L�2ضQ���?�eP�guD*^�n�d
_���sع�^�k�b[��W�Hz�!;Y��!4�f�2Q��c��\!*�>R�_F��0v��#j���~m�}�e�q�go����"׷�w$}�'m2��� �|�d�@��7e�R����q����*���^-�޳�$�vHĈ�u��{��LTS�+c�V���"l|����N*�˅bf"���qv���I �ķ"7�hDo���"�U [�����Ogr�R?�4}<G�&��T��sU��H�qqF�s�nL�08��?1�,u<�u��ϫ�Í�N1A�������_�"�Uk���`�Nx1u�V�	�N��LX�4�S��"�.Q+Ҥ]�cCJ _��H����z�m��u^�ie�u n����*�١���Mʑ�E�c���A��Cl�����	��C�y �H�(�6_�(3X^8�w�L�(�z����w���\�)�3|F ��%@ԗ�[D{d`_i,����ݪ.����K�U(��<ST�� ���P�vcl�U���l��^��ݔ8�����5�
�gtNR�n�ؖ� ^,�DnH�\șY��n��� �~��N��9��$_x���x�>��(��ȋP���$4ڋ�R��n�t���yғ�ڬ��k��{^��S�/���#�=8��S����4����8�:�\�f9y�ȡ����겞\��8K�pC�|q�:_��������\V"eOfH	�fď,27�puS�Q��|�$wʫ{
�m'#d�9��f��O ��8�IXo�^
��6���Ej���%�j#f�e[2��9�����A ���T*{�;]��칽ne&�+m&!n(UZإ�=0:�KK�x�hX��<��\��\�����`>�z$'GA�9���Cs���`s�z���/"���AM��3$Z�*�R�o��P�-��]Ǡ�F+R����>vs����>����_V@Pq��z�o�5�f*E�0�)�t4Y���6_�m`��x���Sm�(�({I)���	v�WF���rÆ��i�����i�U�����^�Z�5����u
��V����?1�������38t�Ow$2CV��߱R�A��o��d��?�;�r �����Y��R�=����A��ЬG>S*�V*Q���N㎁Ό��q�b��p��C	b^�G{ �5��-��b�f�ś㘲���T^:�Yݮ��b�����)z��nD�eo� g�;V��oҥ�7x�yQDG'���5���ո�ػ�L����iX�n4X\Jwl�~ӓ�&F���� ��8��%��b��ͿLm��M�pW�I�X�A*@|khlI�%(w��[��фu���ww�M~Q<bZ{���.ˡ�<��GfX��m������ �L�U��oѭw��Hg��C]X�~��mPg֐F��i>Q#���Fܳ�.e�S9�;������k/�I�AQ�P@DvF�"7����ۡ
�>��y�������c;g�&�M61�xn�~-\�xix&?`����l[�K5Ǐ�@0�C<l���RBf�Ւ�ض��������A�y��ܮ�ɅҠJy�V�$p+��L-}y,�\ě���@��eP*^gY%��k_=�����(D�Ҙ�JK9�`r��[)x:q%�x��a���S�]�;a��Ad��7����kd1.Yi�Y�M���Q�sgM�o&{���gE�=� I��f�d��VS����{���H-R9j͈�g~�W�W��CTE�鮿���:yoaT������Bc?���tf-d@-HrH��HfȖ���_�Y�d�]�G4e���Z�) Ǎ��d��1߂��n3>�/�6��`,mί�g���B����[���>��'����-8����ԡ��6��'��,>�8������V�0}�x�{��o�0p��:N��.Ɣu�XL���8�nӥ�2z�v�I��XEz�tԫ�U�oĮ�9tK�O�[�����ѥ��39��x/�������v�W�+�}����
{�#93l)��=w��K�5�=��'�H���?u� ��o"���|�9{QPw�ą6�	�;�XfS��U�F\�z��y+��@�q��I+��O^p��`�gf
��4[��$�F�O^��Ϧ�#��/��h6V���5i%j_��L�l(@a�;�����O���({�4E�O���5iRA��!;~����-����2���֮N��n[�d
}�i�.D
Wϸ���@q��\�M
��ר+�:%�(�I�����z<��[�#a�4�ǏYHT��F0�K�����Ǩ��U�H���	����y�^@��`}@<o�d�g�ED{�!=�i�K�*>�>g�02)q�d2����<��4u�S���{���q"��
vOk��}��1:���b� I��O����Y�F�k8�.OJe��2�Ol��q&�2<�<Q��3��\�A�2&q�|��#�`�O�|r^��a����a��B���_�v;R9�/7�]EY"Nh���د�F*'���O��|^aA�Z�?�1�'F���H��y��۞�9��r�5y�XKy���{}F��)�0��Q̅��(imOȉ���E��PsWH��`�p�>o�������Ϥ���XC�dCi���_L�2*Z(iw�h��m�Yp�����W���H��*�n��3�t�_�S�tU+M�B�b�/d|��q#�I�F(s���XD�^R'|�h]Yq�̆��2�uO
m3�������h���y�Tc�9
z�蜒�|�3��ǖPI��Kd�{>�^[U�#���y�d	�tK���l�&�Y#��LDDk��}Fв&�p[q��aTxM�Ah��$��5'S0�����5�.6c��zD���n�ﬂ��d�� 6��c����@]#��8���2'~��z
N���i��5a�e�9W�����B�lڗ��%��5�	3<���_�?��i�Sޝ,_0!��RתF��(��<�>*ђm�H(3M�8�
��:X��&�ڟ��<A���[p^k��E'e����0P��e!���:':�r8��,�Gl�7rpϪ�8x���4CV�C!L�xș����q'}b��˓����_BG����vS#�.)�l�����!�Q���"�(>��v��\�!��a���Ʊ�w?�V��ԈB�@}��:O7eCg�Rj�)t��^�9�.m(V3��7;N<`(ʹq�1��*_�Rj4{ �Eav)?�D2�������)���r���"r�Mg2�ЌTɽk���W�P�����:c�C�ΈǤH^�T ��L�b�A�f+N2[�̉�(�g>�LC�}ll1x��X�ψ0��]>����� ��ft�O �����p^���g50`WPz��o����Z8��݊AJ
\������B�r���l�|B�c|7!)O��=]:�s:�'�mF��s�R���[+d4���\EV�����J"��K�����_�)<p_�Sp���@� ���W�� ��r~��1_:,�fI��י�G�U�0�eQ����&SO�-�ʱ����j0����'%���KI����t����#Vj.��"x��jo��ٶW�Ki�3_���.�Å��(a>,3�O�Kq=�� ?��~3�x�	_H��:��|B�I?����Q ��#
�o��p닏UPݤsݎ�&Ջt�I#�w��9�8�=���N��Y��6�9E�����. ����`O�\�Ԍ�����.7s/E������9ܓ���*�'w�=�� a�&���t��B��������v���H�<c�߭iPo���>�/���r� �d�� ���8�Y�ë��8.(��\@��ﻥ��Y��ɜ�E��!�7V�k��(�de�Wƞd
�K�����x��D����.	g��������1�&Sˋ���hsY�Y��W$lP��H�^�kb�_�h?��<T�|���^���T��?�@`K��ӆRzV���$���# >g�lX1EZ���6�"`CC}� X�������Mu��L]���[3K��X�E������:���Q1\�G�哈8�ܳB�}(g���>$�GV�p��~C� �ļռ�T�7ƈ"�^���
0_v$A�-��-��j����J��q!w?z�犣^ڹ����h�
CK�Oʑ1�<�Eݭ��d�.��r*W@��Ƕ��$=\@�y��J��hWi��u˹u�w�F넮�S���X�\�EjQp[��cB��D�q���ŏ��L�&}q"��"�f2WH��� 6yb� ��8l��1���Ez<�Rd
�7�O�r��DKJ��.5���)VS���4M��!�*l�l�T��*	}��
#�}�FC�6ZQBLS��U��qr�f��6���Kj.-U�+DE���Q���� Y>�fl��[�t+OaPL3t�7���D�f���G�8����p�"K�)�/����*��{�er��_��:`���Gw�sص[���IC,�A��ͬp5�᥽ݼ~��t�.�Zڠ}�2	�j�\�0��(vZf�6y^M����8����5uw
gQ:�<
h��N1��!O��+�S;u�VYP�%f�"���e �<�Zq1.��捗�5>��N��ĭU������r�1����1e�M�gq�G$�2���TO̻;�1��o�E��q��Z}ogP�2L5��}Ғ��`�#�i��y>FV[����3[�*��ɔAU%�^��v��#iX~=:�H��	�>�U:8[y��{�ݖ]�yJ>�ˇ^!g�.),:��0l0��n� �o`�>C�y~�����h&.㟜7�Q�66��J�s�����d����^�f���-�}p���(��f��>2}�u���-�ꝕ�ҼIlIjqI�4g��K|���L` �#�1����������J�ڐ�j��9x� 'n�_7��ĩ�{���`�R�^�	�����z��m����������GH&���1]�-?�;?qt�*�Y�gI���+��=�M_.*�ӽ�׀�sy+T31��h��.;����d��ڵ3]1�KPD��Z)�47��zj��iQ�2{���F�*NCI�R�w��Q���e���bFy�ݟi��(��U�U�z�
�ڪ�h^�ƃ��p���A���ʳ3�Q5GP�o���.Q��':���75���0/5F[Ԓ�����8��`��&�+1��F�^�^9��^��	q��2Pb4����MN��}y�AnI��rX�Ϙ�z���q$�:~\�>���F(�
<�/p�����˰��� 4�j�����F�pFWԱ�O��5q�+�NuQs�H.�-���M���UrN�����'Ƀ������7�����M�v����j�T�=y)E���4yG
���~�o\��V�Jj���H$l����'��`��5�\�_�O̇�<�\��>����yC	��x����/_�h7. ���4��#m��R+Gy5����*�i!1/�)��{xz�.�R���=��l*c�p��"��zq�n�,����v�̢7]1z,��fH-�+x�4�M|47&��r�������;�:��xN�®��$O�Q�x��Z�7�9Q��kͬg��B�����L�D��Cm*ׇ���g�gk��q8�j�]K�l�Ķ�\!]b>��Q��@[�/S}�*v�`Nt��VH�_�Y��=7�뀬I{����nCpUV�� $Z6ZU��Nʒ��aF�y����i4�6���wՓ�K�!1*�m6�E��8�oG��#P!�kz�~R����{d��:���;��d�5<�Q�g6�[57A�
y���(�bC�`N��!�~������m5��D>"ђ"��I]E�MG�A���Bf�Ar���9F�����ʞ��Cl��x6�p��G�|�u�ɟ�^R�8ž��3B`g�LI-\�p�D�i��u��>[i�ϵ�U�I�������
�'��_�>үM�0�}��°��ʅJ((�]��C�Xo��涣�����N�F��<�ֵ<J��#}���t�6Ӎ�JCCi���ƃ�
X�5����i��U��c�R��p�����& ȫ��3�Rಃ����TŘĶ�%8�0����.�p�
�P��z��u-N�B#� ��'� �]�t�V'{�J�__޺���)j�Y�Y��B�(�Y��	r>8ѧ�.���S5~e�,D/Q�F:��BH�=FnƧ�.;u���,S,{��G��Wu]�Q�T	�Rw��P�P�~|�T ՚ p��G�u���kk �C=�oT�<k���7|�9c���T9��W�h.v$�����U{cs9�
�	R��Җ�ԌU$���Ϊ�&O�Y����d��4v�XX$��rA���9���@ɫ/,���RN�o�lQM=쒜 "����z���ra�-/k��B��q�&��i�L��Zʩ&���~gR7x�8�,��Cg@d2��n���jr�bÇ���i�6?L.Q$`������']��ӏ>Ԏ%�Q��i��<�O?Q݂b��1��p������	��A#� �ޚC�Օ�<LA���.�piR���9;p&�{��ס�+n$��v�z�4�`'��~��8
�$�Ik�:��H����L3��[̵�_v�������$���M���E�ț������]���I�����I�9�?H��5)f�"���̦��
<�Ӧ�4 ��uy)��N�d�z�G:�m`���㙎���I�+��^Ls��|hR=&>��_[�:M���Qڐ�Ư��F������]x���_��?7��+�J�T�,���7[wG���4�n�=�$�ǳ!�g�����$a_k�Hs~`n�WZ)+,r��l��o�d�� �c�|�%F�o��7i8=aK�X$�o�wʖ�[������9���t�᪶iH)��Gcba�X�K���E��Y+�Q$�]x~ߨ����1�ܹ�׃�=����� �>�4
؎B�A�aVq���}VKrh�,�3�}z�� #v�?v��2r�N��s5r���\�M�!s��R� ���i��~���%�P�����I�/#��Yۑg��p���6H�d&fŁ�Tד���Ir0����]7����XǄx�ڙ5���N��+3P�d�s���{ 5Ar�}$����2�w�H����` Ǒʢ��&����9[
�4_~�-m�'#�5(N����R�â����-�5�r�_��H�Tk<�g�?ٙ�ҭ����)⩓Μ3
�����.:�_�9�������Hv-���� ���	�;�0�=o63j������ �z�@����lt��x�������q��]��5�sM
��[�i�%ȝ��Л�5��2��}�$�k�Gy�I�mz���m��t|�޹�:���<|������@@gP�p�-��x*U��#4��DJ˚t�W�b�����g�oPQ
�1�c��GQ������Ǩ��Q��ZM����<���1�(��,��nһ���T��xy��-��"�n�^fxN����As�zS��b#kq#,l������U�G9���W��(#�Nc�@���;�n]�\����ʸ�o��QΨ�q�od�-	@,8�s��}_�қ���u���i�{6�Gүt���y9Ar��x�W��,3���8��0�h[��F����$+��b�i�n�O��y��3�aҝ�v�C�M�~��ֳ:�
=���b��*ݑ���ªߦ�h_��j�v�)��O|F�/b��1�h�|�n�җCۈ�q���
��d.���z��;����������j)��d�ֵuw�-�FI}(�o�B���ʻ�Ɋ�Y���xN|��uϝn���>W��c���wu�E0�����>��e����>�}[EJ�&�|nEu�����W�r/�1l�;tb��;\�[j\�1ؽd����GZ1F[tUaٕ�{i�=�k ��n��-$�o����f+�S,jM~�M!S�j�q˖B#�Q�ǿ.C�:\��m蜷g�����"�:P�z�a����aKI;�u���׭d"L�(����������28+@������
�������@t�է.�uJ���0���'rkզJ{�����| ���w$����
M�Z3�x$��7]䳮P����lO�Ip7=�����yǕ�r��W�x�^_6O��`H�z����+{Ck�I������p�-�}�}��EqQ7h�Ώ�=���e�ZB&UK����g�hR���5lѰ)�_Y����ۍ���4�^�ǣ� ^2E/E�mǒ�� ��R-��Mq��|	���������qO�!�VȈ�3b���$���':޼����_p����۷c
��%*�Y��*��9�Rz��V�n��_����\�w��_-zQہ�^���HA��>왾(9�18�d��j���(���Ց��C����=R-5�O�����u�N�zrJ�`a�p�M$�Gr��Z���7���ә�&�G�:�QW���B�PRN3���K���V��U�.���v����%���ƣ3�6�����rn� gѾ(ż��VpXY�����̦��-	��'&�O�I@�c΋�|.
�aݰ����tbp�/HYzE*}I�t������=1ق���������:��6�膶b��[��*��e(��v~�K�f�<���ѳn�ӝ�^�0Yч5�ۗ/H�����fÂ����E����]?�W�[Ȫ�]Z�臸:�s5ܳb]+W	+%����������~0��;�P)D��TT���Jٛ��Z���;��Al*�W��Q&���-Nz�4^L�&�;�ڌpV��L�_=���:���w/�tؾ�z��
(d����DC6-8�v�
co!��c����~�~4��
b�Gsۃ��_���b����9�6��۵�P%|<�8�R|��;����\�j���?��%������z����sU���n��Yg�~Qc-e�%�U *)D{e%*�0Fǲ)���+?q GR�#c�+E(���h'�XB,R�n�W�ׁ��&n��H�ؒϫm@��؞��?��g�Kv���UiT�"�G��� k_�СǓ��¤̡��q�Uֺ=M��wOf%k�0�+��M����md��k�V�͈�ʢ�>��TڇΗUm�����]�<D�^�=$�M��&��U�M���[�nx^�$�;LW��Tq�f�@�?��b:�4lnz"���b�¬p���g�o#Ph��2P�ƜY�r7�ʺ��Y�h�C�s�\d�"*P( �^dj���|&S�����˕x9��X�'!����K�TQ�DHb�| r��\�aqb�����$#�w����e�P�@���"	������+Z��C�Ғ�i���j�u�����ٺ���� HhD>%���Cv��&�r��VÚI�TWLJd����j1�rX�hk����=��|�ZR_�ixE3�����Φ��EZ���"A�t�ͷ3Hh{-U���
�7��U�]i�֯��1~<�o�M�N�!����#f�oI?��AAf���.�5���8om��)�B�j�ê}Ʃ��B>�ﲃ���&�l�R�I(���ob4�jC�/�	�ےor c�b�mE���4�a}Ѭ���Lb[�4��+��HΗ5g
�#�
�W��]����"P�+xGS��.��:��F0q;_�*���V�}���T���������Y��)��xB�2B0�2���S�Q��&�`�_"�*}R��(�����O�eA���$�4F<�����P��6H�"V��H��XN�ׯZ���󵜔k��E�k��C����{���Ą����G�J;�7��x��d��2�hq'�[�&{LT��ei �_@-�u?��}�=�K�]H*#�7����@�<�����i�iY�`�����Hdl�Y��FU��0�N,���O���O-h:]O�VMK�z�q�J�i���Ѻ?mRQ�Z��4mzNc�*w�u�6 C:���jܻP��h9!ګM�$!��|�&w�ܧ��J��l�,nP��X&���`I���A�Y�c�C",��G[����S�����m��N#u ҝwj0�ͻ���0>I�e07ǟ&���Ͻ�����"�k�$�%�Ǳ�dۭ��a�gDҲ�P��$g�Co�uȯ+����,�Am״����ןa>�w'��3N��n͔lu��!��=���~�}���!�Kg�"l���w�Y㐌�`�S	�+�/~����q**��H�y:�1��K6෋�mj���w�_ir+�T�}PD9�}�'���q��b2������H�m�xG]ye�V� %�a�P��3vM�x��r[tlmp��'Zu][ {	%��|�	���1&��J=�@��\][:Z�b'�k��r�o�5����}0ZȬ/���Xq<;�1
���#��ܪ_��3�?�wʵ���b9iV���k��k��ʶ���/Ȱy��|f�3;Cu�'���ٮ1����$�r���0;v*r$Ge �+��ҷ4������� @?ra	�K�n�	!��|���Goݬ��q��3N4D`0�hR�i!��S~�@��iò�.�(RX��1���	�{���8Z�&۠$[u.��X|՜b�*iU�9��������Q	��e7K �=F={���~�;��-1�Z��f�;���ݨY�M�j�C�_W_��  �*�@@)^a�Rɢ�'9#*V�%)��F�dT���	6�qK���V1QX��e��kۼ-"`���y~�8c��X��vF�f4?��l���F���E�#����#jr�~��+��م�g�τ��{J9Nak�ZP �KQ=�S�+yʍɫx�E�`�-�,��F:5��r�m}����#OZ�Њ�~��<9��P4�&��Bq� U.�Ss���ְ�3)��zX?2m��co�UF���YG��+�^��̓`���]v��^PPK�_7��!�`��ϙq�U��!.l��6�aU���\{x�`ǂ��.9}.��樭�c5M��X#&|���Ϛj8�dj�B��͡}7P:�{�߻= *L�,
����>P�뱩".:�x��r4):q�[��l�h�i��F�+������!�iR���/="9~����7�9ӚmL��&y��Ӌ�1g��`M��硌v�^�:T�����	��<����䨮z���㭋!��� &�����[-%�gL���OGOэ߈��7X�H
�$Ͽ��@jx��)mw�ʌ�8㈭��3��j���	�k�KPyP�{L�\Ht"ۛ�����"��l�x���9C%c|%�SP�4r � b��&��G���hH���"�	a'��M�"X�@�3�HP;�:�e+�z��;:��E����s\�Z̳�u�I��e:u�� pݘ�g��'ȇ�E���Rs5����E�߹A�q̰�)���F�Ygݳ=B�Y�Ķ7S
�VqX�k�#Ƭ����	ä�/`XEЛ�������~ Y\�V"^�VK4q������.���ü"<~�v��Z�a�!��&.%��u�3f�@4������aQ��*��`��b�*�d��7�.���D)�=�k�N��I6=3�%���qsз�=�/�8����!ה�G��
|Z2���������RH.U�fK�>�OWL�V���D2��5��-1� 3�]B"������F�'TR�ӊ�e��տ��A�h���E�x��'{#�@����?�W�]��@��8���}�t�2\��)�ne�g�����˶��I��w&��Q��Џ+�Q��&��Qp�Vg�E�V��
����:��;��x�����$�jJp��8��tt3�qT7#V���1�I�y��a���;�u�W^�C��Tk<���z��%�p��}�u�(��uLS^E`:���۪�x������ ��ɿc�6�߇^�`�b�V�m����;.�;iߠ��'�,~���م9w��T����D�(R�Pr��a���q��}&$Uo7��t�aCp�vT|�D3�v�|I^h�+�a<��0Ѣ�c$�;�S���Ӟ������S�!��g�BQ��eTp%�_�����3^���O@�-)7��;�_!������J���>����ǐ��Դ��Ʊ�F���2V:B'�S�v�p_bo�a��rP��Ռ/�yO��+��ݵ|�i��KO��S_g�b��
��D��JFΝ����)���<;�u�v�x�,��^���r<��NEμ�10z��d3���^_"P<&�?�#��m�}������!u�9�Ȕ,t��#*LI����[?W0��UX�_g�`�sŖ�y��2Ք�b�[��q|v��G�����X�S�(� 
)��v��=H_ �:'��tˀbu��iM��3��][�N��e�9Q�;0L/)
VH�5U���R��_+�%/_�R̉6� T�IF��/r)&�!�����|�A��:@K9��!(y@�W�O�����,�X4����as��HY�s:��r���x�h �p�^0	�|P�M �YA}�fܩ���G��{vBEφ�U�F�w��J�U��Y��9�u���=_¼ʾ��Xz`��,�����9�R�*���PT(���%��2��)�z8$�x��B2�v����)w�a�]E��(�A!Ϧö�f�:f(=���Ɠ��d����L��nE�#)ꍱIWQ����N���!l7]�/�xQ�����(�cЧ�M
�jg!t��(�_��8$��e2Ԯ�|�^�'uܔ�r��	�M��3���{�5���Q����`@��K �xƿ����pG��1�����xH^��� �Zl��k�O���!+�(�}(D�k�����	�&�$X����*z�6D�L��W�W��K>O�����
��/^�=�;}�@4��n�~j���'�
�RZ"�y(�Թ0�Z��"zȱ(�fl�R��ԗ��#�@�du=4=F�\����S�k4����ՠ;1b��[g�`3�� �
�ڜ�;��ʌ�>e��l�~v����"W&���=�YΩN�\�?~��q��墚�5���2(����״��� #���et�=S���,!9��\�a���L"�ƥ�'ϨQ�eF5�]��]�`��S���AN�6K}$�AAy�.��5��05rvWږ\�B�}ۯ| ��KB�:8N겕�w;e�[ʦ��V80�ɀ����!�k�՟�gZ��v|�xЁ���}K�G� �P	5'k�����#��5R<�i�&S��Q
5���j�m���-�~d�%> ��$d��:�H�*b��di��@?@��҄�c��6(����a���Qf��$�`C��a�|PR�2�Wjk��C�ڳ6맶0��<��uRC����3;&2�I��P���L,�K�.�<7 �W�R����s�T�9:Y�/��Y�Y��߀�# �>�;2"X���Fi=��S�m���8����7��Ӏ�7Ro9�B"}������9�FUטS�8�����2|�=��|@��ĩ��:C��<}��ʵ���r����WN��2ԙB��00�����{�[V������/�d0T����O�G��7�l�i�$����0�h��>]�b�h2��C��&��`�Q���S����?���T��==M֗
>��>G
]��6a��-�wˡ��?1����ꌗz�jy�3V������R4�[)��T�:2�߯�$�	��B�od��YM����n�Dq<5�s��8 �������C�W٦�#88��u����!�7��2�<,SB��)�R��,������@�Ʒ{ι���{<$,J��`�����^�^L�dE�<���A�����9_����h�n���������F���&��¯8E�1�J.�y�v��,)����׌{S���ʬN.�	����5�i!�H�6AJ�ʰ�u<������|�$Hu��1Eߧi�y�7�u�h^���8���2�O+��}��k���t$"�X1��1�����t���)t���9����+o�r�3���Q�����[� ��o�?�Qt�*A�09*�A)��u���)��Tu��1�=iy5��L�X��"�Jw=1��x.�ECe{�e�<����abJ��t�ApZ5�YG~,�a�[�dX����tE��ќ85Y�Z�P�뼋�F�<s�-�Pq��k$D��U�>DR�X��b��4�s��� E��H6�=��Y{8g���� �7*��J��o�A�z����Q�f�"�� cc������f��N���'S�V<��א�l���v���.�h���<1D�@p'�	�
ʅ,��W�%�OT�4�1
��jk��Xkp�Xr >ي�D�2(oV�fO�)6�4AP�3'��|�>�p9���Q0<��~����3��<���Wl��$i�d��' �Y01��3"#��R]��V�:�m\�U�ߵ9���h5-cڨ0�����_`��<S�N�]��;�a��p���?P�z�D�+���� W�ĝ�����r6�F�b@�PwcTg����X����N����Z=�N4�����Q���%d���UV�h݋���a6�f�(��Ks���=H����5���H��A�J-��O�c��������@��Q������V�~�V!mvۻ�p	�W�+sJ�M+�8aH(�٬5�E۹XwȘ3�	�f�����L���VY����mOY���y�=��eV��1l}L�Tx�n$�;Ø�#�X8K�U���˵�(��cݫLu�`���V���E%�K����$�8��7��~E�1�רp-����Y�IY�������?��e
�-�T˸�W\4r	ۋ��P[�G�d�~�f���D��Z�=�4�pȢ�@̼�;�b����9�D�Zn.I�T�q�E�C�����t{}�Do,�[봖\��P.5��TJ��R���<�Z'**�m�;H��WW�f�	� M1��)���������M�h4�κ��\E����ج >�9�O�6H` ~�����l�v#	e��t�����L_�7��8ŕ�3�"�q9)a����
/TR�,�j�ͫm����������u���E��ޕI
�,	��X���d�����[��p�6���%���Y���,A//�(�4�"�b�1u��#�f�{������k���6��6|������&t%��FӖ��@ղI�$��r;]-�+ŕ�>�x}��n�W�E|��ҭ��R��mC(q��D�j�2�C�$�	#��<<�p�8~���Y� +�$�3�f����vϩ���W �߳iˬ3u�xc��|�`X�̈́9Hh�������~H*Fb�<�}u�أ\��)�FJl����|+]O��Zr���n�N�O���f��Ea\r�I�W_d�?��k��n�覈ܔ��SE�g3�>.G����jO�y����h��
�B�q��;Y���4�⤏O� Iq�A��b�07<U<�����0x��l��*�������m�=�oČ�%J׸����8�He���x��k��ȏ.A�zo����a�~r�r���!6a�a�]���΃�QYɞ9�ζŜx�:,M$���!� @F�c���&�нɶ -�!S������Z~��d�ڴ���ޤ$��3٠h_)TF���A�(Ug\/,�`�D�)[�&|�EЌ��,�`��]G��"`hւ�].��e�S��,�z�n͔*`2	e Q*������ n���RT%�Z�X�Z�U��F\�_W]���>/F�"��5�,a75���y���ִ�߆,B%#��W��)��`~s��k�&#�l��k�J'��G���]]Fd�}��A��P��Y��ڍ|�I���MS���QQ�#@0aV �D�dO�]�f��R�%�{|�
�ހ��s����\2V�������v��}-zR�=�ɚ��2NBq���k�x�|�6��B�o��|�����%��Fo����;��1�FV��Y3���k�� ��t�:�+��Nŀf5��6-�u��w�����4n����,@S���P��E�������F͆ɽl���P�j�]���2ǳ�� !Y)��V��* ��xJ;|�jݸ�:�-�ל�K5�pD���r_�#BjM{ڈ�V��JN���Ӥ��	�-�Jo՝/l�r���M_��U��p�o���i�e�k�l?�~�Ơ�w��6l,���^���B^�Zd���P�?(�K�ߒ��w���C�a���D��%���</+��f�\»}(w�@�M':/$J�0D�Yi�C�1��l�VK������jlrP��z��.�����HZ�Be�f���|�fC˱����ya������{��3���i%��@[�����	������	p�-�H]�n��w=C�a��G���bj�I�!�����j r����~_k}��rɲ�J?w��~�`e.���m�@V�
�1&8Zq}2��}��g�ͩ}��K�w�8zRv�z�l�	�^ބ�S�0}��}{�v�$�ǰ��8�'��K�3~�|(.'�l� k!�"O<h�:�/y~�o�d@y<x^)S�%{�h(�y/�G�8��Mc3��9}�{B���c���Ɍ8�����C9�8��.�^��E˔��_�*i�f�>6��)P�ff����Vߟ�#��m̙l�\~�AMi���ӎ�#��TO��S}.�D���J�^|�-�4Z��Di�����;����d��Xn>��+��ԢVk��q\=�֔`G��f{�ƻz^��T1�P�v�uۛ^C�s����ʭq^TΕP&�R����$דj�ZH֬���S�*X�sOMLѝv�R�D����L�&&����i�s� ^�ؔv���t��j�k����O �P����$v��T`H���ʯ���BϜk��tT+k#�����î0�1����19^WT*P���[˞���='ˉय़ �ˏH�{O/�`On�0�L��
�RP����$�2�b@~����O�$öq�@�%H���m���%_��qH_�HZD�f��) {�]#�v �vL?���o�0�&ĳ��|�0P��*��_�:��ݱsD�NY��a�0A��g��\��%s[������ I$l�v|�A΄���3�MP>�&<�zk z@DXvג7�~����=o�e��Ï>o8Дβ�����ǖ'Vx������|�����������j�`���Y��E�w���e���G��$;��j���)xB7%[�3�^**s��M2�s<�X�ά��������r��,���/��%d'p��<<�k5��4|j���@lq�N!�?L��^i�0Ia1s���%*���ׅ2�}��/�dE�l;f���R��#��K�w�}j����)O긂ůI��-�ݵ���"* �2�8��(7Cvt#�^���e�=�Vd���*b>��;�?J�]�B_�O�������o��.�"2i'����\�&s2�2�A����Y筕/`%<ڟPg��)�	q��_�zw��f��/�!=���h:̮����kM��9�n�flS�)������ę��}�HZ|4��2	�6��7' ��%��^(���t��D`.�wo1bݹ]��;���B�W���6���@O9g�;E�K��H���zL��,��
[��n+!VA)Psr����ʻ����t�����Tlf��ĉ7m�'�t�֘@O��t��G�=�K)V�.�f׵î���S(��c� ?C?�v������<����B?i�i�r����w�c��1Ƶ�sq#3x����iҸ�N�dt#���rg���������Ѹv�*%��Z����I�q|������};�q��-�����H�Na���(�'�r��Af�MQaМd��?a`$����Bv�Y��(|��ˈ�(���4�e��y3� �$)����������Iz��\�
���X ���=%�LVX��@�:=tg��Cٝ\�÷gaj�\�jG��]�tN��Gbt�j������g��j@��0 ����|(cd�_��-�q��c�'�-�11s a���~��O�3�Y��6�2
-�/S����#��QD��;��ħ��m�gonD؆�M�j~z����2g��;7����
�(�A��h5NO� *���(�^�?$�s�B�}�3�B���?n?�Oщ���3���>Q���K�ZYh�<��R���֤�����Q��L�-���O0�}KK��W!z��%%����#~ {�7@��w�/6���G�:������"LJ�a��k��׵z��ʁ��=����Kl[|LX#5��#6��-Y��fĎ��WzA8�������V��o�����)%r,u�-w�;F���+_�R�3��C�,�j��,��1iI�h�� ��oF*l�"���!�$�i<���ԙ�+k��k/Z�@|�	������DN
��󐇙����3}�t0�K�>�m�=���Ք՘�M��YG�uA�"7�r�1pw���A�G?��
[Y��
��W�!ud��Μ�)�ӿa��h ���N��KV'xʼ:�ȉG�qn����ٖ�C��!�1��Y�p���a}�nΨ��GF�!Гd?H�61�ۦ6�Fb�^xz> "�~7n�ͥ�W��AvXԡSV�F���H`}3����<���+���Qc��]�F��淰o+J�`!xR~&�0��ƍ��	���o*��Lꧼ脞w��vEQ�](���1w7P��.���=2Ӕ#�����I\��P��f��BrTݽ��DQ���ty�i�F:��\jD���wv�(X�S��"�?�=�ɹs3��*����aƷ`#��-�P��n��Jig{1����\?�8Ϝa��Xˋ���Y1�J���� �T�Be���`jf��~}�¨�+2c>�+��Wh�'�k�/��o��X�7�p+4�IH��mq�޶� m�sA�{�m:��������U?8�u�B4	��_܌���I��7A������%.QGaiY�/X�ţ�t����1���B|;C<��gW�be�I�\4�N��>O6bb�)�����_�N�
�4Gm�>�R��-��]|p�/����* ��t*��k��%�R7m�Qx4D�l��v����@U�h)lu$��5��S�~�5
�W��[�88�Ql��g������~���W"'��]��̔灢Cf�-���Q�ȶ;�4\���#&�f`�@�w�1(춄����n (I;j�[�,�l�L����֪�=��
e
]�&����R���.}9����r�B(����3� �!���G�i;W���3|F݇8��٩�+*�l�Pn
@ٺV$��n**;v�Q���(���7a��CQ�.ɠT�Y20!�G��ܯw��-��'<z#����-ֳY�<nѯ̪�2UWēh��ʩ��:���Բ%ʇ�o�1�az��h1��G��#hE���Geo���OLd��{>Mߧ�ўzvy�9J��a�N�u���e.�~�'m��p�Gv�Q�n�V��q���7�H�1sU��th�7|�w!Y��n�ó0q�����qj�8<f#��CYO
���W����!d�>N���x�ъ���%{���.�C�h_"�m����ϙ�;�{Mu��cD�'��>�'�����2�!4�øQ-�|��&�p���'�r��~sc�W;G�I�|x�C�������*���+,���҄�2�B���У�8� z
k���V�x�va�m���C�Jo������hEQ�=pm��?�yM�Y_�=�VH�MD]�|���m��$�wXv�)>uvt���w�>�\��
�J�@\�y�:��_n���D/�#I��٫y�j`Y��c�sM<�g��ً�\ �x���x�rD��(�)}�� ���=�I��aGXT���T�su�.�Ԋ ���
1nl.�)(1a��j#n��Eh�J�a�&8�c�����Z�S�tD�e�NĸS��WRXf���|�a��>Z�P�߾�|�lłRa@Oj��"J]c�q��hЦg��M�Q��?uI����[�w
"S�+~+�$eΑ��#�e"����] �f�an�U�~���������2K(��R7���}x�^��u ������s1�5�X�N.�?X0ѿ^�_µ�os ��6g�^��aI��r`D���[��%����2�@z9���ƾ#���v�I*�($i�?��yv�P�ٗw<ޅ  0�w�&z��DU8_�.,�5�����	L�M���O8�o"��}��I6�X��֛�q����`I��5)���Wr���L���M��|��e-ބLU/ê\�"݉�M����:�挷��
�����0��48�w�#�@�aQz:�D�Y����6x���!���J~��JP�ͥ�9A�k��=%����z�*��*��:�	�,t���8�Omy����u	f�[?%�0��$������3D��O>�6{p�)�Q�
��ꃠ�c�݆E�(����u/	��D�,ӻ�84���g,���gk��cg4�a͡��*{TL�!����S��xU�C�}�F[�k*x1�1�_GQ��\k�z����r��Z52��/"��`�e�f��̖�Ln�_�	d��<��4ϣXx��&i4�#��p,�~���E"R]�i���4!�J���-a��Ɇ���c�I4�ш���j��i����(��@�����ڍV)�����m;PC��@�����؞\&`�'��Yᴨ��9إ��<j!ݘ�k4��
��Dv$�*E�����7�4��Q/D�	#<=s|��ݿ�jz)�����Q6�:HZ�G���C�L��������_ۭ����SM;���3FW��2p3���������O����}#�+̈�ќ��(��g��g� p��qn�<w߸(�֔1U�m��j�̓O5�(m#��x�>�2��Bo��a�os�������+��{��!M(�E���w�R5̨�bRv�ܳ�S��ĕ�@�lޗ8ܠ�ǖ�СZ�f8F9z���L�(�_(��'{��P�5I������_*٦<9�b��(��80(ig~�ٟ˧��ވ. (���8���vF�8�\`^[�2xkT��}��dft$B�?�#`_�1(��m�
���/�W�9(�+SF�D� H}�G�8����k Y2,n~Q�Ϧu����|��:�t�š`�:k��G����2=������Tq�yI'��x�T�ex�(��j�����o��w$,���,C��f�`�֯Ӧ<��Gc�Ὺ4<F=��M�w�cB�P�2�G2�@�ӵ���m��D+���|5���̿��
#<?.��Pw��<9O���W<�����W��a�0Ǫ���ш�u�DR˻�UVܸZVb��B.|�a��D�N�����AL E#Z���
�Q�����|j#����>r�;0�q��X/^�a�p�	4S�����];�Ֆ��:��;V�3IP��~��s���ì�^8��n�8)�OdfM�:l�v�M�cf�r���7l]���<��B��K.2V5/c&�g�$b �����9{��6�Nԯ�Az�1x��Ÿ��m���	�_	�k��*:�,�SW�s�v[$�Z�S��t9�}�5��i����7���/:Y$��;�(�o}l�f��B5-�p�J��̓�5��a�P�}b$��7�d���tsyn���R{�n�R&m� ����ǫ�_"��g!Q���%�\cZ[���O�Ƨ�pʙ�>�ͥ�wk�7X�zj�/*_h�m��D�a����)�t�X-W�FZ��A�8���,n� �VD�~��j���*��?Ub��X��k$�$�99YT�9y�c����V��t��
��Sc�|6�.^$G)�{��
�nU0��oȳ���jl��;��^����u-ø�������V�m��������8�a�Z�,�I���UQ�� Q���Z�6��k��Z���Z�-nd�����/N
y7?�PG3?5~����0�ԯ8&��ks�������������x�ۿz!��#o�{��
瘯"�N��۽*�{��:4z;��V�#i?��1��*jP�x�2	b��:�Եq�8��ށL2�K<D�p���%g�E[l��(�_�:'�Cr!�����J���m��~��/��0�Ki�)]UN�8/��+��,G �*y��Ҋ�XK�.kTg�+6�G4^��"�,��*׆�1��?�� ?��؇@�.���G���jt0 "b(���x�aC|��ڭ{ё��@�J�CEȫ]�G�A�bcu������^N�|?�,���6	��fB�ۂyD���4~:%,�,�E�͜E`�I����Wr%`Q"t7��r*�!H��^��V-viz\v/������Z�m�21;$3W�R��ƀ���si�Vϭ%	VOٞ�ؤ�X�B���d�h���c��@�|[B��7�$�Ï�/p}�����<A�>����U�:>;jC��TS���x@f��'K/y"��Z�2[=����0�)KVM�}�<XP|�jA��}�[Os�.ߣb�ڒ_Og̳�G�DR�f��?���~�����b9����,@��8����~�~K�_Aܵ��?��=�v����&���ϑ�'��8�#n���}��ڢ�q���vt��!�aϣ�f� �~�^mE��a톡AkG蛊%����� 8ʰ%�ो⦛xOw����x��Sˬ��+1efm̸-y$���1թ��P�wX!�i��ׇg~�W�p�S5�~�*��'I�\;i>�:����3@.�$��p5b.��q��{���o��D8��O���ɾy�����Gߞ��A�ָ�+i��;hZ!���R�]���F �\aи�L�+E܅B�D� {+�_3- t��e��!�P!mj����� FΫ`FJ�e�|ucm��u��L�)\_������|e�¸��lT��e�vF�U�Mrq�(����KJ�[�Qi���g�#=7]�u#uj�f{PP�`Ju�L��=��tH<;ϛav�y���E���|�D>\�����ص1`��G�3/G�����&�O������I6ky�ɸ~�l�{^Y����E�O` F��s%14c�?j*[��nc�խ�6V��?�C
h�> �>�+=^I��d�]P�=��ۖk�β(�Z�-i�'$/]`���˦�a��q��u�)7�����1�Z�{o�Yq����M����h�2�eo!+?�)�]��DUӾ*�=�S!up{3gAS7�}����V�����6�2�Fr�P���y�_�g-7��n�V��蝓�V�k=$��Q���v�����a�r҄��A|WY^!�ۅ������%=�cCT_���D8�Y�N���8�w�o�M*/��#HpXH�I���:����:J� g����T�l����bmD�G���vV��<-�̵�F�w$��Jr�:!�����1vZ�|D�l� �ß��*w�BȂ����	��X����K�R>3�j�Ҟ}���rb���!Ʀy���_t�$�.�-�Ќ�x�	��|;
s�U���� �!��RS� �fʞ�-�y���)K̋�9��������S���R/r��\5��QTR-�~�&3a�g���ەS����/��O�X`���r*R��! ��J�?"��.rzP�l2z�S��L�š:j��vK�2��ŝ����gA��-�}8j���'�E�*r%�V�� �($���2b�%���Hff�bT=������X9� �M����Uo���0}5���p:
e���ٛ�8�N��6Њ`��Ƹ4�TX�{�  q|��^��vd�C�+���Zҙ2P���'"�����x���f��X&�&̕�*.6����/a,Ly+[Ύ�m��H1'�n}�F��6�ڟ�h�
R�����j�^t-��8�7��N̝�G�i|�DP�q�lO<Ϗ���K��{�b_U*�Y)5�ryT�i��S|��@e#s �2�7n���i.�K��/�u�/[,��A�n�ĞA���Rgx/ǳϞ�'SO�z/�%��AI�s�NTE���X����@ecB�ꎎ��3=\y�X�@��!���˷�O�ּl�KIǷ�eٓ��q!�THVH��md]���O�~��R�0���L8�T��BiEqg�I
i�������֌&��J�܀!^��ԒƥςGyb�$�N��	�k��/����D�	��Ə��w\U�>�#xJ��8[*"����`<yi���OM�6f!s�y�n_�Z�0"���9X�>W[�Z��QJ �(���}rw��~/>(X#1���P��ѝu���->x��)�؆!�v��6����-ڼ�8n�� ���k}�*~ܱN�^��~սg[��F��6U���f֍P�nO���&+��!N �UT�\*�&C)4ꅅH�[	�+ưs�d�����CcoϚ�ڗ�F��Q�>}w�y�C�wF�{��"�˓�˽��53��121�Y��6Y�O������a^�(Yl� ��[���m,'(���篵hP��0�[a7��Z�	)p��,M:'䢈v4^=|���'�����R}��9�45���M�G�ʜ��F�7�V,���3��'���B@����E�Q�PI��8��ORAmY�bj�?��H�Sڈ���9���$�Ȁ��(A��"A�)R���豌�mE-!_�'��(�9X��t�9����İE��-��Y���1�F8��!~@��`C� �K���j/N#�B�������,�+��/lm("�j��j�?d����Gy��U>���:�o~�g\�����qPF��::��)�^s�Hg]!c�F(�J4j�]���W*ޙ��S��C����� �S)�_eu�Í0��]l��C�4}˻���o`UT2���rP[����AX:� M0�����z�� �f�y	{�8�����TPo]3$w{w�ߪ=�V���{��A;X
TU(��+Nb��6^�"��W~��y����*N̝>=�-$�����H=������,9q�|� �SM�q�{���O%l_�k�Y�c9v�GR�pB~	c��6�"�p�<[����D�4t�nB�$�Y������_�R �U�W�x
>H�@�̉�"���$��sX�f^���B$<'�bS���_{M�U�)"ϐ*���b�T��70�c���,�V�� *�nk��YV�<�0��HY9�;��Y�@��\�
3��9nu�}g��Rjpum�C?3�k<��R$�@���m-M���+��%f��7	d�`*��^�e��oWy����c9ާwX7�_D�O��S�"���G����w8!��Gű���2�7�1ܐ�\�a�c���uc�|")XN:�.n�;����<���vƳ@� 
]Q�E�������[S�r[j��!�hc�GD�a��T,'�9L�'0'˲g�OWʛ$�6Ғ�_Q^.)�`ܮ�z�֧�J�@��"�]rUJv��D��o፰�f���$n�5�WŞҾU?�3(����خ��Hx�@+�0g϶�Qà�t��|��{W� ���Ë7��m>�|��4:���]Q�-��Л�`�]R��{l��� ��{����>�@�h@L��ZKk�.���uI$BR��vFI��Ʊh�a�܃d�)bF��$�$�S���f`8NT��M�L�!O���9	�1zb}���G�Ou�l�<?����Q��O0O?�U����(a����y.�y|}#ݒ3�#�0
2�����ȵ�1�>y�vUN���`�"�,���Y�U+H��#�#CvRJ�6dLh�����Å(4jK�gS =�s��U�JF �='�*��/���Q�d.��r�O�WnXvؚt�W�d ��K(?@
戢�W�>6xI���!�R��	� �N>�@_om��~fG3h�"Q�At�*�ݑ��E�
x��L�i.T_trh��r����k��(ڨ>��l60%hL�؝�����8t��w�����W����Cټ�1뷅�&Pvd��[BwαW�Ff������n�x�8�2�p< ��|��$�c$�s�F�����)N��a�����)�?�z��_��GY%E�˘7;���F��LV��JG�y_C���ر��W&����k���������H%�� ��Փ��D<�C|T��ďג$�h_����P��=#C_���5����)�5�|�n�s}N.�u� \�q�I�1M,��sG�,G8;��3���@צ�"Q�w����8����e-2xuJVәv௜�ӂ����.�^I\!���v��$�z�*?7-��;�M��|Lp(溍�Pv[@��D2R��qm�ƚ<��v�I��<!�#���*,2���`Zu�� �����Ⱦ6�5�@�y*u��� ��)6�����X)��ԡ�XD��J6����e��X��)����V@�\�H���+�i��op&�	P�����Tzv?5�a��OO��)��|>䰇x��D�$��jt[og�1Ѫ~۴�_x	�j�¼U����B��K=���3>/!w�����4������2�v�����p�"�L=��w�A�J������}$B(Y�W�u��*w�T0p�y���.L7l��S��r�v�2W\f�&�Z�$[%����M1����h)���+3��wOc�=�B�M=�g��-�F��Xb�	b%��bXo�d�����0�u�[���p�،�N.�/���lx3�᪎��o�	�9�2���d|ƥm�P���{}d�ĺJC#�Ϛ�0�A�$�1n$7SR-�C��;q�a��l0�'�PiSR�J�~�;<���
Lwu+��Z�?��2I��>Gk��NZ�,�_(e�*j��|��'������Hِ֦1K����8	�P���	���r�~��۬�����$�9���v{����~?}d�\�B��Á:&a��r-�u���y�l�B̭"�I�҅���UJs:�`�/7��1�Xy.K��ty}�9��G���Ǩ���hu��*�Ʈ�z^�x�o=�LA�ҁ� o��<Z��0v'��t��uHJU ��EU��t�Ċ�xu����'�pMPc}Yy K��[��_p�����Fp+-�A	�W���i��YT�M�X.W*;/���2�n�B����"�B�)j;��rG�������u�������0F��I,.�B]�w b�#L�&Vv�Q(B�b�1�zz��^a�J��8I��)�\5\y�ڪQ �����%�I���ͣ�`�L��Vs�u�FJa��Iq𗌖��/�r���ےQ��m�5k�ج�]�q;���G	Ocՠ��~����d��d��]4����aϖMf:�����NȂ���%���/L.Wm��7D�,ӏ���
Y��Ǒ��U0�Fd��&=�/<�'v�w����ht?:��DX�N�*훭�G��ah��\���y�gz�Nb�-_St����&s̞J7!�S��rNhS���vs�A�����ɒ��~s�zf[p��w \$3�>�Y��cR.'O){S�!Gߠ%�"�l��'C��H��Nj~>�o��q�a���գ�&rH* ?�4�WCr2�j�Ⱥb�A�5��mW(5TF�>/!���{b�4#��HP�!T'ylX��T�˰�/�*���5��µl�}�2��r�[�cq��ڇ�t�
Ye��>�A=����c����tl��s�Ev��"�`�S7����9����Ev��:�mkBD,A9�K�~��\��}�ߍ�#�Qm���@.���1��O��;ŷ�����q\�d��6&��+�vέ|�E_9��q1~�4���f��v�|p��h�!0£j/OX�}mntO(��;՝���#N��UXCr��T�xlb��q)Ш�u��֧���'�.DO��?�W\�6�.�R�Dwԟ՝6�����`�r5�p��0X˪	X7b�Rv�ڢF+�"}y5���2Y�Ra��l�y�S�Fa��'�ɐ^9L,L��D�������A�xC�fkM$��dȃ$���l"����{Ab�諕�h��uXY�<6�{���t�D�r���/moӤ���w(oҮ���&L�_��LYG
���ԉ�R&Ţ����L��~�]Ѡ@䵥F�Z�����+�z`ԍ�	�PRز���%�Z����t����O���N"�`�@�Ϟ�Sy��X�k�o��q ����r}�w�'�9s��k�.���q��qEF~ *γO�/Z�h��T@�!�|�����6V�\\���׌��؞K>uM�K0�� efȢ�[>=���7<�Xt�"�����ݖ\���	>��~�ѓ��������]�q�[-��6+�I��s]�?d��(4Ɂ�ni��S����Gg�QM��8G���'<��o�����]�Q�A�|ՖT#x����Tq�Sw2���e���|G��ѷ�F��� ��m�-�#	?������%k��ҳ�bwMh䵵5Q��W���O��}3$��'��%N�!S���VD�k r�g:.�V�s2Sq�,)����)�BPo�	H���~tjd$9��F-r?Mv�6_"Ƿ��`��ű���竚!��ݐ����	>b#e?u:=�ׇ��>���Nc�� ns�K>��Ī�ǿX�,{�LS�]�@���[�u�m�ʄ]�H6i}��j�G�V��k�은�n�W��C�7�;n��$�mv]�Q�#9�\.cK�>��H_ [�� ��I�BH_�Pv�ƍ�\��h�G=���/�;��f� y�;Kr�@������'�X�H�B��0{s��3�?w�5��"Os���w�������LfjB�����&�'C�z�GT1��	��K� ӗٜ�*�=��J�Αo.�WA;0 �y��?���Ј�a#;��%s�� �M	�P/ܵ'A�J�.É���0�Qb�W�Nl��n���w�����;4�a����L*�6+��=�)Y{1ה�q�#WK�K�{�(���-�B܋H�=M����-�r�xH��ݵZS%��I�@�ճ�Hy�f�"�O�O==bxT�u���
��q_4�$�Ȋ>�����YsǱ?��B����>���0����L��3���a7�����bI�ΒcC�ht���G�>ҁ�B��s�v�l�&���?F�R�S�I�g�j�5ṳ� �w=~����?ʧ��
8&�2K��=@m��M��*B,����L\h١�l�0�5U�q������v�����P�q�OJ#I��f��Ԏ��y;�:�*-�\�$�t)��M���^���Öt�"� SH/9�|��=-��0vi*�z���}̘�ŝ�dj-�X��*%U�}6�j��|� }o�NMՉC��p���ǣB�30#� ׃Γ>�s��>Ļ�"Ƴ��q�����|]~�QS�x�d�u��M��]џ����e���|x�<�-86Gn���O\���i7����%��M�7��_qP��d6����i���tR�.���$���c*��,�G�5A���!1@h/hG��cBE��|e
 [�|\�w��*a��H��WK�!�Nq�&vR���	3]��(µŇS��o��fN�w*kɤu�e�j�~��1�NU(���:�]��W�z���.On��?*���7��Iȕ�hO%�������A`���hEv2�*��G0��'�ro�w:N�c[�*�9X�Hٸ=�!{�x���$���Л�:�(��,��B��6�/��(yo����i��͸�~!����g'����4'VD��Fd��>_����&Wcڰ��{�����,���c��M�==�oǛ��7���K�5g?>м�t�NZ��h)&�y
�NV���"�p�O�yHUft����_@K�пDi|b"�dS7�lъ	�'�������4B��_@Nt��o۟�B�!�i�<H/"4x5�ѨoY�E-A82d
syR����4��r��:�E�WoQF]s"��\j�y��������ݝ�Bs���zjzb�J )~�M�F��25_���7��&�RC��o%#�m����#�����,��h��G��lV�O�b�ۛY�S�<�b9���j�֌�B�D�?��~��A�f�����'�,��y%� 7_��RH��-� ,A22��S8���O|\;��(�Xp��R�n'>+f��w8?���hf�������x1�d�!����EV����P�����.;��sU+��ij����bh�t�m��GVp4i��]F�5�����4#�~��y}&��@���/���Xcd�֙��g#q�<R�ǰ��% �E��ao���N�
a�rrq3?�
B������HT5'�6��}��c���#�jH�;�2�5�vc��=\�z��J�R�s�o}{�b�����ޘ.��MU�,��܉5�<�j�%��LO�����]���ئ*M�;_<�k�MY�N%r�Oa�/S�ۖ�Ǹ[� �$���z�n�2%����"�DCU�g�����?�<o���F��?��w�*«����;�q���3kY8��&{ʎ�,M�Xu-�e�飚�va�HKeVҺT���؋b`��g�AW0&Do>��;X���}?"ڕ��
�J�;χ����O���Bd�!-�7@�o�E�]��P��~��9���ޭ��Bxd���e��V�$�p��MĆd��e�F�ǁ�Η�U(i̲|[�`j�+�lfn���^L#�*��j$�E�`b���V��y<����{�A��y�sK�����䊓��v��#���r>��~�9> �+n�?�����]!Ca�6j�����zE�ғ)r]� h1[N�s2O(��8Q������`�m��9�Hk�m��t���IV�8Udd��cD׏.�R�U������ϑ�s�AN��ˢ�~Z��5-Y;����u
4�Hwn�D���J-
$;O���&��.��N!�0`k!Ԡ������Ym��o ����g.5��tK�ٍ�i�ԩY���jA��DES�E���C���e���ȨvD̯�,{�9����$�{s����bB���_��y�Hts7���G��ݖs�ǐ����TU�*�l"x%�^�U4[�e< [��1mu��n���4���~����I(d��ڧ�5 G.��)�bk���xuVn-K��nb���؂
�[+��B�%�@Rӥ8�뷨H��jWl
wD�Բ�����nE�D<m�r���NSZ��DD����[f����74��9�{*\���ح[4!���m��	M�EE��)c��h�(�ip~\mܬIAI�*CWs�Z��jw�	�f�s��r2�dУ���q��KH�	⑇@�9���,�?�r���c�۽W�w9��R�{*S_����H	&�Uh����B�@��-�m��WW<���f�FŃ��%�K�@��w��Ɓ�xaB(eO���W������_z��Pl�헠�:��]�F8nRJ؂�A����Eՙ�mC���D5Z���X��J�R�p�=5(��rB	Y.�Yl��)���4��(��z�c�'쨤amB$ӳ�A��֊<�����^)E�<-E3�|T�� 
���S��O˺�*�,��-ǎ2���	�q��=�r�]h��yD�M�F�..�K�B�&��9���o���0O��m���"Vo�n�kZ����R�#�E� �e����<�\���R�dյ��ݰ����9L���b1��c!mn���ޭ�a0�qz7[<0Ȧ��Lhw���4��ɵu�M�7��W�_6;c8�5H�(�x,��}X Ԙ�2�����C�1���,������S���� �ف�iؔ��z���z1�%�����s#<@��F��>�����kz����BF�T�F�	�F�M���K�W9�1tE�`y��ba���1��!�tG��%ek���9�y"Z'���Mx��t�4?�����y��EE�H��R'�;TT������Htb�#��H�R�8<+8�d|��wz�n�>�.J�?PW�'j�Ƣ�@�}��{SM�WO�n���L���bA��U�3ڝ�p�#��I6���郴��R��~��-��V���a�~��&1�$�2u�~��,���� ��1�h����Q�n� }���W��c&�Gg0��V��cM�3���,RUC�A�����+�{(�>@�q:���3T�3F�dG�8��Wx��C�Zjz6E'4�Ůtuk���(oE�Ƕ�gf�"r�U��.j�`����V�=xQ#q+�����/�Z�H��]?�3>U��J�w��9c�Nΐ�h�U�G&jIw��21�@�Kd�ט�VKP*,Vn�6i��͆��wQ��\�@��2�a�����.bf�,��������W�~P+��fOݹ�62)�a���P�{$]������̫`ED4}zx��
���2�G�(�l[ �*e����Uo�&i;�K��@,�I�b�#�&���P
�^:6��.I����	0+]:��Kp��)@!��/����]l�Ij��d������(��q�˴���耐���dq^�Xvƫ&u�ӛ��|fά*�o�6{�gZ��?- ��,����A@,#Į�4��iC�Y���O/���3<�j�<̙�{���,�t�gܴ�/yO[r)Q%!������u2j�`���$���L��ҫ�B"0Jc���R���}�Y�=��A6�&�<y�H��-��s�Os�B�
���\�/Q�	���!ѿ��L�)e��;R�q�C\���U���z!uf�o��_څ�_m�@���ƃ�W��P�nۦqq��� Q��ڪj����=4�����/�~ޱ�Oa?ޕ������h�VA��	_��,,WE�YEӞ�t�?4� ���8�2P/��h��h��g�	� ��Re��5R��^���'�cV�����nK!���I���.��&��"_�T�F�7�©@##i`��np�t��Nd�ћ���n%����@�iǾ��
���ѫxcג z:=q�E\xA�(�j�ڄ 6��Q>Xj�2��Y�m+\#�bE�E~��Aí��Y����/\7 h�ᷟJ�� �#ro(^�s -`��Z��f��:Ŭ��{�}ӱ+H�����\4Č@ZI��]������q��4��~/�qC�����[lc��M�� �$����TѪ���*t\��r�Zե�X[��1:�n��f�s�?�2y��+"���i�O�Y���J�T<�;G#n[�;N�P���o2�r(އ��5�)����ԯ!��9b�V�R�3�q�6xq1aO}=R(�vs��'����F�����f�4�$D���t�x#�YX62l�V�*�n#�+�b1����:����q�k�}]F&��,w�1
�{}�L�̒�u�t�
��Mϸ�i�(�<Q�+���;�)�hi��!;'��Qs�6������	�/f瓜�L��l�w���9eAʗ�����D^��y9<���e���v��������!":�g�03'k'b��f�i��M.���0�+u�I�Df`�N$2��a-%	��,S���8��T�� ~��V��4n{HmN6�\�f�>>Z݂�>x�1��Ȣ4GeՕ�� �Rh���k��*A���G�h�������tz�΂���~�6�斨��v�Y
���{8L\5��Y����/�>t�G�VWq�N+�h����e]Sc�aÂ-,ڔ���l��a�	RNĆٟ���
�u���f[�Y���r�N1�j� �Y�w]�]�b����J!$v����k��4�q�K����YA�%P�!�b(e<�(��� @�4�_km���@��lŬ}N���e�XH��p^*'�t��oj������Όҗ�q��5S�s�k��{)F�� Ů���x��iH�u@f��K(����*���,��%��k{�&=�i�����nl��j0b)��)Z*�J�*���E�3y������*B��� Չ�C��y�7[D*Pv�6��ɯ8��Ks�yxD���WF�0.d�^�lA��o��`o�P���Ǌy��/�,QCt��Њ��/.��$K��k�do�87eGեBa����k��G
���H���ۉ�X*�+�)�H�>�����e7� #���ٞ7f�M�Z>����ꍊ�Jw����E}�q���?S��9�Oz���x3����gO�jL�S���~\T�ɷ`bEo�Zb0z���8_BB3Yy(�uJ���i�y����XE��E.�nN߽�-�NCg�D�F{;ߩ��;��v�Vn�c��@�wK@�|�K��G��O7������.��>��c�<�젺M^�=7�'r��tu������\�OD�������~�[Q��kїp�b~u�ic�"=0��(x���*���*J�p-W	��Q|eo.O�o�U�a�O6�!��׋Gc�ư[u��2���)Z��"�3 ��q��G�EZ2�I�8�*O�i� ^�`1�zt�H,�9�vjA�D[y�!̽Ō�����U47h�GQ�zP�S�l	ϒP@�T�Վ�S��:=�����}�S�u�)>�����nf޺�:��ARP��6k��!aն�x��F�8_wjN���im�����c�
`{����[��!���2�w�M����w?vQAJQ�'|H΁��/KO���<�
��N�Q�����wt�#Us4T�*�^N$��ka&}6u�r��_κI�70��$m�_s�������������iD��#��� "M���'0ں(��9�O򀞣������ef�?�9IY�޹UKA��Bj�=���Q�3�Y}O�`$�&�nF��{�`ud�add���1�V^e�0����?�	��cs�V�X�g��J�������Ŕ��k���i>������/%���7�Sb\W����l��F�ߢ-�Y�rH��?]ϑg<�_�+_�;<����;��-�a��}�$u����YK��=S��"���dʑ�-�K�)���P�����>��I�TBv�j�u �^�������.F7`���J��o^����VI�)y�S�^'Ix�`�ݍ��ܙ�����۴��#�����鮒��8J�lY�����q]��ǩ>E�7�O�3�[O�e�I7���(i�h�u����,ݾS�a�.#NM�ر�\ �+�r}	}\�~r̢
\�)���]d��SH���_�l�G� _z���O�hbY=�J̶����R$����<��%�+o�Y ֑�4�����T}����Y�h>��0��e���-���ӓ
7/��F�*�0چ��g^��ĮP��jk����
�w�m�ұ���oBٯOnf~[t�]�l_58%7 q�ujU�qkj�&�DUc�_۟�fe�(4jI�놮޿��QN���KL�GAl��|f���/^�]TM	���^�U,���xn��Je�~,^�qɬd�f��d"�1�E���,x��(���
;����#S���6��2ͱ�.'�c�r�Rz�����(�,�#C
�f�.q�zgA�.����<�P�8��nܚ��"��8�y!�I���9��iY�uL E���0���Y�dPa��h1PT�#c����$+��	�^Ϭ�/^�e�$�(�L���u;r=�����|�����]���7�23:�W4ڠ�i��I|�DsS�U�XE帬l��~�+��6t=�u��Qm���B�P���P�j��x�wB/��H�=b��.�$2�Edv��d�h3c.��ƣl*��!*����[�����~�DB=�8�c��&R%o�>Ɔ����pYɒʔhP<<���ĵ���p��i�=���nq��<��4�E��ym}b�-!�m��$��y!� N���
JH!<��k0K�{�ޯ�O��g��N���"�݅��'Tq\����0V��0���cMҞ4�F�D�ӵI13�=��}nY�����,ㅱf'V٣3�C���r,�@�Zn*�x�����(c�~zN/���h��3SOL$��Mz�F�Nxkt-��j��@��iϚ���zsՏ��j+����Z�5%�GY'Я���!�������|�l�r�M��彑�M!�IE07�T�0j^&��}�U2��6�,��[�TD��I�Ֆ�K�<a(�eĢ�B�#`����Pv%=h|FC�h~.�0\��*D�@��9�d�נ�\><�k���]����V(���,���@�����
���@��5����o$�c�ԩ��ڧj�~���*�a^0�]�y��>,J���ĩ���<Q������7?f&Ť �"���0�њ¦4SQ�+�|(;����L�zﲞD�R�6R�D��I)�d!Q9�����*�=����b��Fr���J�!���&��7ln�
�u�KU�y�=�:����9!N	h\�2�&ZY>K��O����}2�|�c�@����x�Bj��r�a���StS�ͪb-�l��.타�I����]��b;���Bt#��ߴ� ���X�n�����7F?��pdLX�ע��]�D�̇g�P��X����7�2n)�����Uv���|�=w��[;���Z�G��)��Rb�[��Bf+h>ؖ�C�|�"���-ʖ�)���T��Wf�����.��*FV9�{P|��t�;�������$w�+lk����Q���"T�����h��~�J4[?l�|[<�T	8S�|cc6�,���>��u�h���B��p0�Oh��*Y����$��-����m��u�M�Y�1��&������na	���f�d����d��ޯqz1��5w����'��&�D���V����-mo�Ao&�X�n�ʡ��v��e`�Q8&�z����Y�k�8&j#4��h2:��Y�7#��8�0��Bo���g���71HCʺ��#�8�F���\���G3�Iʠ滔�Z軶��˞�������E7=$m_��B�a�i4�"c���|���"�M��r`;N~yᮭ��s�	�P�-}�՞0=��/�\�k
E�J���1
�ܤUP}��F��+&��Z|q��j+���НoP�E�qt�(M��o���o�7�_�4��]���\��ٯ��XX���;�	�'W�@p�� �m՝��$0�uHC��1�`Ӂ��F��r����	��]�������d���t"����	�!�Sh�!�sF?�����0�cq��L �G�F�?����?P�� �V���]�����ٜ����4(7P��IL���q}�^��^�j��/&T<��-�����7�i���F<z^+�� �"G�Մ�<߁�����C�}XZ���tE�r�9�e�Jn�&N;���đ�s�&�#��È���ei:�Z����CW��?/H���X���x]��Ĥ�ՙ����Qx�\~�� ��]tm�����!���OJ0ȄH{���K�l�(;)?�7�������� $1�C'���7�0R�"���~��:���z��A�-�q6��]4:пK�V}�2���Mݺ�`��(�PD��?)�hME�((����~�<�S\���NA�����a{�4�h�0�j,Wf�� �K痷������i�nU�A�^ L��AW'2�	o#�G!,��pb���X��R>V�m�&��/�(�>|�:��&�H�+�ot�A�\e)�����y�w�X�3�8<F$Ƹt���Y7�^�	��"S��S <�ߚ���UjR2˪8�y<'G�$�������_��Q��ט���늰����o@���=VN��Dv����A�E�˺����c�Cg/�:��N|���7Hh�7J�!m*���F���oŁu��Ȭ`Q�V>��!�{z�ſc�W�J�k��>ק�Ta�7�IY�3�D �Mb&ʩ�ɓ�Z+➤�叿f�R��G��
S�P���[t��/���Y�s�̦Z�h����!#��hF��ǔ��̨���$*�v�X�Rx-��}�Gn͓.�~���!��"�>���*�g���T��4�,�Gp8���gz��/�)ƫ���ה��j�ͦM�5}O�ȸ��{^w��Ab�Z�v��J���	s�=� �,��� S~�2�Xp:4�j�_���x�I/�D�k��O�4}]"�����t��	�ȷ��n{ ؕ �:�&�ɛI��EN��T§.��ur���,ΰ��&x�&�̆�:K�N�����x�JCf�99ђm���?�w��:CJŶ����;��MRx�}�N0b<��_��-N��GV��&j���Dr�j=s����O���=��DY/v������?\�qxp���촲���9��[�H�5�Z2;}���D�;�6$o@;Qi/��4}B�����7iF8�҈݁���t1X4�h���r��}~iB �pgqv�w�&���Ҩ�H��(a8 W��n]�ؤ�0�ދ�K�`A��X����(�3��/n<�	�O� 5���7��/��Tj��0di3�ܤTe�c��Qu��9ǑP1�4o|Ih�J�f��,.9yx P=-?%�G��)�p�8GOt��5�	�E�v���*�P�>�ˀ�42L�o�z�hPK�	�-8@�e$�������=�F����>�@��	-в��t��o(�~�����'�)�~~G^�s����"`1f��"��6R7J>0�=�Le(r����-�5�s"��lo�â��.�ԍ��/�<���~�x�K����$g�tm{���`�Lv� ��Vܺ�����\鼣C�,��{3�飙8�i��v���X��,��} �Z8���m����x;��=��C�\ϧjjy�r��9��fH���6yգ��o�����	�7�}��cՄ�����Z�tfC+��fq��0�D.w���>�����>j��3��L�ynT��+��qf��L�� ڗ-[d���0�u������p}|�w9�h������M� �%���v�i)`90٫������ߍ^ծ�|JN���G�ޠ��vօWQ��cǾ�v�j:��T#ұB�$�? vԕ�)�
xC��8OT�#+�Er����E)��mh����a�ڤ�Şp�o����c%%�K֍�Kg�B
�+�����_�,��F�7��3�
z'�o���A�!!�ת���	����NW�k��?9�y�߹�b���va�r�K��G3~��]��Nr,#�?�L�64�Jث+<pǣk�m��*�a�HL����|i�%�����>#�U
0y�ĥ�z;�ǁ{ŝ��SV��& �*'{��E&1Y��>���?��B)�t�U:��o�����9��d-允�aR�_�t��ǈahx`T�,�g����ՒrY*'�v��<fOQ{�y� &u��O��5
4.�!��q���<��]���>��V?f���/N�zz���#J�ᢄ���P�O��$��:�^&C��Xh�S|/�4ؿ��sW�j��C����U�����@H����oa�����=f��֛,���#\[4���[�,t���YBQ����MH����0� �5/ ��|�٪�!��R�!n�e��E�u:�8��r�V�@�Q��
���E�+�7�G$t���y��}*ӷ䒠ƯW�t'ٴ|�@���H�4���)��D*W3�b��R�GV7}��u���jx�Ƒ&�7V��5���v&8[�����u���mc��㣅��ԏ#�(3���[PK�o�4������oM��;AѢ��I��-0�����Q�*
���L�\hR���)�wy�9��E���h,y"%�H���=���w��]p�||kJ�Am�\���;���b���\��+V�k�Hp�S��vn��?����e$�AI}t9jo�3�����5?�J��/N�<�!���'�h��$�L��x��W���k�r�X1M�:��LQG����DF^�x�𳟳��Q��;�����GD*[aO���"c�'�F~M�����h���AF�����z!bZ%w	,^��z+��@H@2Gگű@#'S�T����l���Q#���G\��gom�+d��u�$^?�]QJ9�55��OHf�|Z)Y��#L�އ�qI7�ˢ�Y�Ut�n�w�[F�z��ğxz�� ���[�9��#�m�/����0,,yL%�`�QS�s ���1�>�v�8�<��4��ٴ?z�����Tv�{���]�-U8�w2��_���݀j���
)�̲T��=�+������"�DKG}QY��ͥ��<ys�#0�$���@{����)Dk�tiv�s�P�Q
�@�Y�7UH��Wy(��	����d�ϓ���M�"��(�fǙ<�a�u8+�2��A�(r(�u�Gp�C�*�{�>��}ɯ��[��~*��ꜧ&����e,� � ���J�Xd,+��dXf«�T{����똟�-���I{~F�	釓o������;8�iV��}'��υ��ce�:�}�<MF�)o��3T�$pʥ �9����.�/��:��Q��"ω�Zf�n����J�M��_��S!q3�s-��i_�l~!�3��;k���KV��!jg��̩Kj�����ߺJ��p��bC�9䨺%��p���te4|��c�'a||U�<����K���|L���"}-M�����Ӌ.��=*�|[�"! 	P��!��^�>|���.,���l�}�`oS���6E��%l�Y�А���S��{�@���|��Bp ����Rn)�x�)��fiX6����aeg�V�ݱB�ǬJ���S��<#j�0G2b�a~)��5�����5GSH��Rb���$�eJC�ԁɧt%�sCd���Z��{,������%ՏY)��b���$Ms_� j!�o_u���HO1x��4;TJ��]�b�� z:��@�eLT���2�U����k�p���.�{7	�T�]���d��;�3Iv�6����w�	� ��l�,%�kְP~�)&����1��@S����)Qq�{F$@�He�@;�g�\?ʅ������0�vǷ�b����Gԭ�@��`,W�:���;���e�[�N���.��޿)sVc��
��'�އ�c Z'��k��ŋ�X��h�T���8�����o�4����0
�/5�XQ�Gw�p�F�6�
�U&	�O���e5�q{!�_0��x�V	��SS-�,���6k.����B^2x�%���x!�ؿm��#��7b�`e��!:�N�R5XA��"X��v&���w!���[�s��x�)�J@�\k$S�J<�W -H��RS��
��O�~�C��O�فQ"Q�)�,�ϩҌ)�q��</��j�z�Er�aWm5$y��'��k`��dC^�R�aHD����<�fh�w}?����=�&>树C:�B�w��Q��I��lk>bsi�`�J\�k:v�ګp���,�����+���=&�5�<��]�l��8������<(���}{KT�niI@�%hrnW+�e����h�K@�,U����
���~������H6bb�a&���g�-"���4_����b��
v�u�=�8��N�t�Ed%����/��7Z��c��L�/��6/Y$���&e6��$Bw�x�Ak��O�K��6�7i+�!Q
-�(ӼM�t��k-6����\���9�N�zM\�nĆ@������`��e7E_K�{@b�q�YD�{0�N��O*\!Xl:ܜ���w�������2+�B�����N�>�H��2�P�%
^�0^�m�����`��1�n�{N�w�@7?��	�3)F}\�F�
8��V����Q[�k#��Tz*vx�H7D��A�CR�|r������
��8I�M�t��a�[����Y�Չ�ZrA@���O�X���:!��ŃG�<2^����Y��H�ؘ��Pv^�P���o��I��\ᙨ�A:�h�b I�7�
��������e�����?�Mۑ��?Og�lI�&�|:S��u.��	r�Rf��� ��E�+�ߔ�� ���ݟgʈ�D۪��Z�m�d�-�HI`{.��Kn�����SA"c{�m����k��M���H�v�g��A9�O�]������2d��i�GjL]��ś���#�a�E
?�ky��B&�W�4�D��DWǘ�D *A�0:m ���ϭ. S,�x�GThU�
��Bp#H�}���anP�A���a�X������s9f(�d^��Ǚ��B������tyR���!�$��`��3��%����20��5X��FV+w�6
�(Ă��}�2�F�֌w�71�N�K�;��(�3�Tzp��tFqK��Gډ���W��>T]�Z��} rg^��ʏ�+��@{�^�3����?�A���q���ËK�U/�}d��������-��u\ص�8�$�r��zo�A���:K��z@�Å�$O�`\���#7�\��%��t�`�����M��󭮄�����*r&>:�gX�XI	���Ś�٩1�w=��}#��46N�A��q�ց�X��/D��,xeչ��9M��ȃQ�Tѹ�6(��M��O����>�FAc�V�nA�lU!T���*?����CNy�/��R���W�O
���������2z��bF�
�z�'g��4�5��;+A����R$V������_�}X���tŅ��<(/���݆6;�ν5��G_�	/	W�R�\�	��QP���d���B�F���7͖�@�{�D����M�9y�w��R��_��1u���|zEY��yR�;ыO#};�9L(�1�ư�[E�-�Â���%��a��S!��<��jk�q�~�4�5�PG��%$�[E�bCe[�mɋ3��� �oS�$ڑ��*M�
�L�c�q�rw\*����y�O��uu{1���E��`��V�1��Ly9]��[Cq��l$�[���c��C�P�t�|���̝Ps�a5��L3�*�j?�e@��lĞϛ�vE��d!9��EYRn�(;;����LKޡY�RbC�2����/Ʃ!�NR�O94��Ap-AV�0, ��7�(u�	��å�0{�
 �v%�ҧ҈���d�6X��y��| D"���UK�Z��>�6�����ٜw=��U�RcX�Y�A��._��"�&���dX�h;��Dd<m;��M���K�+����QK�^�5`*�"��}Gr�hװ�|�B_�x6l�^�AFL�m5�����}o����%�X$J����)οrM?q(֢t�����eG�|Ɓ^`D~zAN/Jh�엱N=���ġ�="z��Π��M��A�OY�{Q�����?7!8����������_�����?�	�)[f�.]d�#5��_���o\��b�	��F�QC��y��i0�?��?�ByZ��G��%Z�Vjw�t����(uٸ�]Dk���q�2,{�G%8�K�D���K�����gUsd���^�Pյ� ���R�X�kǇ��$R�3��LO������#s��D�o�eaB��0�L'>�S��R��ϖk������W���;��/ >c|b۸B� ja�p����Ν�W���`EE��0АG�'��%7��'MG���݃�h��X�-�z����F��d�`l�<(#��G�+��J�Ѣ��;���=���þ��R5�b����"����&��s¬S7��������F�������j��x��$�8Î$��*����rƥ�yI-g�Hx�%�?�ڴş �'=�!'6t�� �o�a���S�͒=Ma�R>�ul�ۈ��c�O�S�C;$�ҁ��%���I�MW0u��!���)�'G��4{Z��7�P|T�jE�E^�4�0%�2��>���
qy��V�`B7�������5_����EhK�v�t��컑0��f:��%f����;1wf���״�.^s2���u�/>��4
��P�[F�K�oj��js����	
�y�R���h{�>���'f2L��Փ�Qx-����y(hѠ8�~t��6��a�n{�����,��ww���Re�h}���<�\���LmB�B��G`�"�a`s�o!9���4E��R��}CAKQ.ƀ�T��R����<(X.�Q�i��_1*[�ec�Vk�!r��ȿ_c�k��<�DJ���C�A2a�}��h9���L��?����Rݻ�]�,���3l[��q�O�KU�;x-��#�hT�߮G���T��}�-ϳ�wjgA�A�9t}}LS����W�%
�0�-w�ߠ<
�o��I�^M�	�z�n�&3�����n� ��+�G�K��b)�>�69,�S.}��3� w�.�x��5&�0�L�� ;�l=BF�PAo����	k���V'�5��ۤ�S������9�����=֛��q���^��'��,���&�+L��D%#��y W����4�6�b�[|�$reD���D�oI�c�raZ�TF �� �o��U;�m0�:���O|�W)�H���{����-P����;_�8yn�����X��9_~*�V]ei孀T���Awx:Ѥ �˗�
b�$��)�/n��G�BM��q��p�v/Irh��!��+^}I��h�ҵ�fhRN׭y���j8�Z��F4�6�O��'�Oh�y����6,C�ڄk�&'S|@�c�����K�ߞ���/�m�Z�}gH�D��QV�I�w=5���ƣ��3(�m��:7u�I	LP�$a�%`�XZ�yGX��PX�Tu���&���!���b����[n:��u�#�$�$���x�;O�J��i�R�x�a�ѵ���-���-����"�`Rc(�~ɔ��/���f������d�ˣ�)�	�AճZ�>���S4�,���:�XEu���CwQ�ERX�x݃� #y9_o4�)�F�-�8'G��ŏ�ZP�6\Y��?*�ꈎ�$��*r�N�8�QGM,VT8�����ts8^=��o~�
O���3d�4\C(�y��-�J",˭�j�2��u�+fE���'���[�����{vD��̔�����eD���uY!�h��?�,I���͂����ſ����%~�!m͑�okɆo�*��)�]N�ؠ|���4*�(��ܲW�p�K���Zr594V���w�g�#{�J��
⍓X�6��N@Z�έ�S[z��;���,�[jO����7���
�T>�h:y���fҠ��Iތ��95Z�m��D��_���pW��������F�}3���K�sL��6�y�4�C�!�xPD�(���Ŧ�������"u�Q���.���*4g�)6�$K���b��^o��je�?c�Ja�H�	ˎ�1�ނ��8L����l�f������m3y{2@y~�Ӑ?fP�vd�t�)�Y��K
DD�,�AKsM���}	vW�wC:-����@T��梪�E�ʹ��`�.>�ճ�h�Tv�V<����Z��{h�Tm��cDt�8�>�nh���h;��^���	��>ܩ�����(��T��x,���_z���7ʾ���^g9q*��}����s]J��`���0�P�vz�J�p�DG��7�ś��u���⟞�g�@�a��K��I�>g��ef�����w�lS�c
�g44�X�f�=g�@P�YI5�����'���E��"�9hZEZ-GDU�-;MBȟ喿�����l�ߖ���Q��K��<���H��X?g9�,G��#ؑ�^��I��vj:���ݭ1�������D���g��C����e�n���·�!�yIO�-�!"��q����S�&2Q,���
I%�,�`7[|���-T�GH�u�	����5�l�yJFm%4:d��勃��r������v2(S�FV/s-�$���4��%�1#vmö�H\�8����Fe�����t��p�$�r�t*8��&��q�HtE5���-l�t�{����ʹ���q�ba���!YG9hm�+���*��7I�W���({�Cd�/O|2��e��E툰r�l»:�lZn/[L�d/� �俉~��4Ol���ƥ��*fZ�=JQ	Q��,�D��RA�~]b��'`���ɋ$�\[�D�b�� ��P!8{���y��ƪ�:3C����������xikXG��?s`��H���F����wD6 8�P6�>e]�c�F�k�lKے��EAТM
��Nb�����2��7mk7������	���g
�&���	\-�v=����/�:^�usC�����Р���U��?uu)��]�E���k�q_���T��4�Y�^�����u=dnrZp�Y�d�|sV�z�uڐy�{7 ��@�_���ݷ]�^��1\����@2��y�|���՜$���4�v�G`��
�N�:p�u��"�7�R�f�c����D��X��*L=�3&�JVW�E�.��ë��%bLEV1�����X�K�Y���	|��w����Jo3�� �xr*�>�}8�eD� ����uW2��k�zv�H��u����7O��P
��U��ޢ��f��
��*!.�K����坟�=L?>x �j���=a{���U��}�_;<���W����ȷBS:��5�ߑ+8�d�+��A	�O�o��p��c�I�O9�p�`��@��3y|�'˳\�^1����ll뤳��I�Am��4��� �n��`�"�!W��������S����J�qeg�1;�>���>5���(���9�v����C��� P��5 =� N�� �-5�+k�}�tR���C�0`{ߗ���"F^{B|r�Y�3� ���z���Q7+�Ì�(�c\A�օw_�9�3�u�x�ۚ���v��sh$�� �Ɣ��P�17��p�!�%�
�o���ߜzG�wz��"�gf�	�CMUx�
%�X��\Xz,K�����:��:��}��:E~�N7��e��h4��e�Sg�I2`K~�?��P;��y4t��d�������K��P���P��Dt̟�E���߽�l�DA���}���2D�!5����H�*;r�c? �ȣ�-�G��0����"�3��Z�n�gv��B����&���f����\��Yt�"p��M�e9b$&����P���8"gsף�]��GrK�[�_�Dǃ+���]�k�ˈF�
5�I�b�ê��k�ܼ�h�VS4O�$�r�h�Ety1��)J1pm�'Y��=�w�Fښ�eU����
`���H��JZS������R]0���.�.�Ƙ�9g���~�p;	���'r���;t(�h�1���0��`�S]��"� p�[���f*�Jo Ӫ�1~�5	@��:���fT��GX>L�!����g�b�dYq_�|6�+9���f��˴G<�\�X|R�t�h=�)F	m����G�����Y�{���*G�@��+P�X�"S���f
��v���ߎ
�L$�d�NϤb���g�l��FKjUWQU~j��y��g����o�݈h!���U&��-Dt73g9~����X[Z�9$x"Q��73!�>{]���,�����4�1�V�|ռE!�����Gee�R����㽌�X��TK�&Iϰ����ݟ3��(��?��1����p7�-o� ��1p_��_��d���˝w�������O
!�N캼�̜b�dTV�����w͔O������qDq�C/ch�$�H�N;�L7@����p��y��uT�;��F���ܭ����D��bOr��k���o4��"�:���<�l>���	�������3�^.؄��34��K`�b�d����ª�`D�H�������h�2ҫ�+<��7�P�e��5�)�����5>0�.�k�7��.��7�|�6Bۓ�#��t�����d%����M5��ϻz��;j�o����,|S��{�nZnk�����嶖�����D
���Z��6��~P���u| �;�R���G�p�=I�F�����>"��6v:%u\߼b���H�ƣ��E�o����O�O��C��U_���ƛ
�m� '@ e�4��H>��b�� �'m-N_�2A1V��b(��)2�Z(�r���
�C���@lζ`�Rnӷ���ִ�9��4�Ȑ"E���.7��{DA+���,	�!��V�1�T)��(}k��
Q�6�Ȁ���x%�]ZFY���	
W@C�f����Nn��]�J��m�}�g����VY�C &��b���^��YE,�c�,�4l� �[��~�z���N�6��b�v����ᓓ�\N=�����)\<����Wv�g�'�TM�$� R�$Ά��l�������H����T��f��d��J��!#�z��в���g���MXt�=J��b6����?��~��c��-J0qEx=�����͎m��:K���b����y����H����H!Q����B���q>�Fq�����A4W:�r ݳ)�x�c~���y��N�T�{�(!`Py��J�m���_�������Mb��1�
�?q}�ܯ'��JnP�G'$�FU����(�=�j���lI�I���p� �rO+n��+�duɖݳ�܉օ[�k1j��l��*y�ު��yo�����~���vd�{H�!���#��h�*�l�/5�7 �vF��шF�V0I����e}-F�b�����e��d_��!KIE[}�jSia��<Ñ�C�"gG�K\��C��Y����Q�=ps�Tü\J�'�F���ۦ��,W�\:.�t 
�i(e@�eI!#�׌ܨ���+��I:����So����HK���h�p��X-��R�!}oCrd��:!@����M%Τ(HbqyT�b�����9��H��[�R�Ì���Ѭ?6R��'�H�z��X�Ikl�?e�M0%�H����ؐEfw��ÊEŉIk�j�@�1����B����+�];�'Q�+Pk�����K�������83O�j��}`��!���KА�:������'m���̊���<��|�ة��׼Lf46%>�E;�X܇*�=�vt����U����ӹ��ű�,�$;퐷=�㷈��{���b���Z�9!�� tN'�^�O;̛�F(���q�|�".3Yn؍nݙ�
!$�jwk��<�Rr�#[�1�i��@1�����.�~��*�5M(s��O��_D�'̢K�����hs�8��=~�+`{0݌�t��c���ц����l ��BP��?�������m�z�Td�mb���1	���ʽ�}��c�f+fQ���[���&��<Bdoy"���x0��> �)na���6<��������RLg�ZE"k'��P�@a �*�5p��{���������G�䞤�s��x��a�v�x�o�U6Ou�Ɏ4�f�t�8Ư1]���6]�ᐹy`����Z��Br�q��.��^��aV�>��+'x�8_��ωWa�e��o�k����U�&6��N�KN��C��2�"���c������׍���8u��U]�z���0�P��5��~�P�͡��fQ>�ܯ0�0��5��R/>��`���k��C����H�����@D<UGh��!�^g,�T^�U[�h��,���,�ܡ�9�4�Ag&�{3At.���Hb���%�-K���(:��Vs"�k]�l��{1���]`4��;�%�+&����[����Gk�-$��s�)���>Q��=}/c[D;1-A���	���,���R��s�ͨ����Sidn�
1�I�mڌ�����k��O�<��үL�F��7T�����ߕ�����Q���O�ѐ:y���C��#kz��	����V�»;�>��aϊ�nK��:L�Q��:�N�#�?'��~�w���Yyh��`�OZ�Yb4�3��=�޸�H��-�������YNk�V�HCfB�9.~�č�eK�/\5P�c��7���iZ ��%+�����)ɶ��8I:�ڜ�ݥ�@�Ы+di��+�Ȍ��W�}��=<�l�_���,B[�[7�,��4��؜���o^\+��f�Lΰ �{�(�_A�8��6 ==%��I{XY,S�B{�㒒2���a���g#�z�z�UTᤐ�,G�]w�{�(mZ,����{�����eHd�k�[���ח	b���2�r�g���7�N�=��n�3�&�L��4֥���}_5�?�F�A�a�t�e�=w,�X�fڔ���fV��A^<}�	\�_��ª�9�M�/�xxh�'��E�_}N�֒�R�k<Ea8Ȅ�Qz`��f��������UL�r�#����CI�g�IO��j�\
��j�k7��'���**fħU[;1�tzɂ!����M?(˓)�����WEA�=E{Q������Z^���3z+o�݅��F:�ĉ_��y��z��>��O�?�W�ҒA�2�1N��3� Jؼ�%f��f�����/���p�`�N��!���Q� �`�Ǎ &�Tݬ>!�ȗ�tPٷ���1j%1�W���ނ�;(����0� `�(^�uS�Wpox
s�?�����{�ݕV4&��5�',�P�p�u�먛�gv�����P��d�i,���l�q�s���E�(���2��SQ�~R�-�Ȉ�;���]`"��Wj�Լ~/�'�X�-���T.�=!{�����W�0�j�܉�ϋ��qS`��[��Je[�����nX�_k��x�>�=���nٸ�a������_v7��?A�З;Q�]�?���̌>��>�C3��{ i��L��l�ɥ�EqP~;�YjI�b�{��y�&��!�tH�i��y��JC�.	�FJ97��)�*��BgkV�L���.}hg�P"Si�9}�ܯ��+���~,l�y��xs���7s��~�T!�6��B
 �v�|զ�zlbx�w�:���
ҷ6���@r�� ��,��n��J�:H�X����@�qY`>�R//�e:�����m��]_���^�,���&�ǀ�6f��BOG߷��W���H�_�[S�]߯G+�:0��wղޓ���:��q���$I�QBz�8O[{�&��Y�#f�.�a����n����ц�`�A��Q�뽘��~����al≒��.Վ��8� ��-e8T��Ld-K
99����}����f�7O�����θ�֪�u��v���n&�XdB���Q�%W�-� ��{�f< l�;��Z�8BO�H�&f�Fˎ�	�!y
���L��q8��M�41�h�!U]���mB��tL�g��%?9AS�큐�CtO�������ْ�7ix&�Vت?C�d����B�x/�0��`s�9�J��3x=��%� 2�kq�������M����I=�.5�#4^g����2���L;*��G��O��M�;�.H	s�"����WLZ�T��j���Dk�q��b&�΄�Ơ+v>�땎5��.G)��u�j���Ф�YѸ��n�]��_���x�dҭ�5c9���6�������ykG���\gF%I�5B}t5���=P�gT8�m���{Bp��M4�h���8�}P�f� c& �B G����R�J��R�xf���T��_��LW6%�����Dіd�#}��m�"� �+��y��3ʈ���ׅ6�n���5j�������a��?صnXEWU3B÷�D:�Ĕ\�s����3���n�����aŜ�p͑����%�T�3A!�u`����ک9�_�ƍ��Xr�	�J$�G����D���"/���Z���e��x�RSMMi12hwp���)d�~\����o�`�\�M��^o[9C�k^��6�y�O���W���V�N4�_�q� ��,l�{U�N=6��9����"mxrG]ߜ���Pf�Mf��{=飶�v����+�#���3'jѤ����o١�e9��x��$)����:�q/���ԯ�y$�j��DD�b����c^���nXG6���Z�8>�\p�"qZ}����kl`Bp�f�4����]��I=�-鎹��}�\f����`r�W]ŎƟe�Vx�M����7�g&Z����t��-�s�362/N��dך�R}����b�U�W��օ���x�����GG���r�i���[ʢ��UY���}��P���4�|�<؅��_��="�0�n���V�|	�$bw"��O@6�x*,[ܪ��1fj��g��i�~hR,�V����~	,hx�%�b���u�^H�{�!)��P�O��ftH����'X.��蚳�
U5�����@���F�4�&�Eez��DZZ�n�>�*�\$FK�*ɿ��Fe��.���[õ1�tҵLg!�Kx�a̼�(�UX��Fw��0�0�Ɵ�Z��v2�ж�N�b�9���
��"'�N��
{��>i��k��y�sU�)hkL�a�כ�Xt�b
ir+J�E�F��Oh��������D�b�G�%gS*�X��&��:y����;,��YMq���׃^8a�OM0{Ǹk����i�o�w��
&�1���\��!�����d������E�t��%O�g�Z7������u<��>�UqΡ'Ĉ����j�#2�ֹr�z�>�DO�����AQ�f8�I�ڌW��m+H����'�fV���&�g�g`�����{}^#c`����l��?3���J��\�ނ����$&��m�*&G�~mM���h*��'�!�-۫��\K�&i��=p�/if`���U"`��<.q�I`�6�U�k�9K���N���cbXU�ڳŮ �GNPk2*�Z�r_4�\-�A7�cG��(*1
К�#�O�O��$Q�2�"�Yѷ+Eg���G�ߐ���MT��*L:��nFօzC@��0�1��u��I����L� 6�Z_�%$�[S#85).qclB05D��@Q�K���m�d�(#��H���x
7�Xɫ�d�!��0�&W�^͏��a��q&,b(ek���	��0>�]PM��
<���B��M��s�R�_V�I7�y��(�`�VD���_�����Ѥ"�C�!���K0}ɪx���{l�4:����z

aV/>�b��6�WәV���+k�C]y3�����H��8�.���(MW��;w��2��Fs���L3<r�X)x\6]|��Y0����!��H�J�#��W���t�=�|��*/Dq+]Ba���ʝ�|�� ��zEѹ�������S��r�,7z�����iZM�K���sP���|�
��p̍恱V� m�q�8b�	��7.&"��<��`��C�FHq�f�Ԥ?,��	mI��m�V��wz���S�Q���{��	�.\���T��zf'UPt���� X��>����P��������=ԼzKЁ�@�{�����х�y����4	B	���;n0�Syn��z74�\׳v��呖�D8�$Z�*K_V͕�d 
��!{�x�~�p�$��Laa��w���O�^�Śݘ��+�k���s�*(&M���/�O /�C?����u��!i����V��"D�E�S���U��&
�+�K��L�B��R.d�y�ksz:�і������e�i�uNA�����\x�c`%v�rW1�5O�qn��8�>\(���))��*qSR#���=NN���'�ʪ�X����
d]!�����` 㟽�K�)5�$�l�	@�I,7GfD+o�n��8�j���&�׃J��knz��z�M��岲�~�����j��!�beO��j�0�~��l��o�-��uj\_��O�Im��3��4M$`��(k���@ڿ�K�iH���"�f�P��ɛt�&cM�=CzJKGC�3r�ɥ�+M/E��9u�9�Ps*�k%����9A��;�j*�'�7Y�?M��C�:�3������k\Kޟ��lj�u&/�Q�=?#
�_xX�X� _s��鿍,[@(*��C6y_C8��2��e�%�
%��)�]�M$
n�8���u�%a�MT]��"�����O�(��H��)�y��U�a�!<x9L�����ݢ���]!qm�B3�4��J�B�w���T>�E�jgӖ�H�W��!���˒�M���۴z�VN�u�6��{t���l|�;"��. �=�	�75�簼�:L>�
����mRUk�H*$�7�BU?f�v���4��g��Ư0� ,����hޣ�1�����`��&���B���D��/ݩ��O̖`Eݱ]��0�TycL�W��	��.��� }=���� �:�x �/jy=��϶&�%�J?"�lk����D�|˲�X�F�h[1M���[hZ�5��h��Na�N�Z�>Iׂ%��w��7Ы��/m!�J%%q�I�Q(�p�t���J���Q@�yCچ6]Oa����o�U=�2 G����`�~-�-@8�]<�sx��%���E���9��s\����;�{��fa'@)O���|��XT��b��P�*�
��&�!�:ѻ�|%�'��j�BNC�`�/Ѿh��tA�c�WT� ls�u;ۙM��n!ɹ~�.��گn�ķ�ņ�~ns��N�3�ev";�Ͽ�s�m�+���³�f^��;v�ߖF"H� �r�T��u�������������;��8(L���5��p��V�:��8���a���0��َGs���^ޱ�g�`�/��e���I0$���p/cU=;�~�K�� 3
=�B�����M68U�����'��2��Qo���JP4��)���)�s��qY8��<���b{�/��p��dA)��}ϟ����.�4Ƣ!�8����#B�}��	@Ag�����uB3�zVAx��2����.��Y�Jjx�x��S��U��=��Z�a�y��|r#IV_dQL0�h��c- M'�g�ݕ�T�@$�^AsASS����+��]3m�e��2��ԯ{�?�ӄOQ��3�)�#�k|I����L�?�6��k�[̰S���A�[-/��9s.3�%Qw��X#�ceD��	�b#.h���������ia{�6�ma#����P���� �(I4�@�	���8�Jb�NM��=�ϓ+�@���+��B�lH&��G|C������0B��=���+�8�}7����t[:���3Ʀh�sO��L��iu0�����\~�f%XE�+��Z����o�Nr�%�f틂YFB�ZB&Ã��+Y?�&��<�\���,��(�v�_�#s���b����{��v��0SM-9�B�@�Q�<򖯋�)�aM���ꔯ��e�(�ӆ��p��>V�Ԇ7)��is�B!�.uj1���A@KtШ���TR�g�H����?�T{IE U��U�CuU���V@s{�;�yQ��a��3�:$+�^扼��:%E���V�UO�Fs&N9���[���<O2T�7��A�B����)E,����?z��8��� s��ݯs��5��zL�2xJJ6h��|��Gb�n&�<`P7�_$?�'�SU��Ϙs��doQe-����e�
>���//NzeK�c�<��z��(�]aG�$��
�|��Ǎ�~�Sd��'��o���;A�
��Y�%8<m���d�d�d��Sr&��\'�Ege���<�5�MF��ߊ�X��<�Ӗ���7�ʟ�Ԧ�og*XVv������	">�6oI���.|�bxD_{�?��ݩ��f	*nC�M��02��.�����^wɁ
�;�3��K��a���k~n�}�f�O%<P������ H�2T�9P�/wU����T͉�=��7m*R�
"�/g!�'d�T.�Ʋ�8m�a�4�S+(lEKD����F���]�X�FlG-"(��
�4�)�6�	Q�d���Q_~�*b.#,k�U�U��?G��=��$)�s���ǯz�Z�#��&te4������{�U���wg�E4�x���T���8��ֺ�AW���R�״ʂv�ą�]���oT�!O
m̈́�=q�d�r�'"=�t�Y$�Y�8��u�ǹM�[^�1��-ɸ	���@�.�^2EZ
h��¨�*̨V��񛣋��j�$�>g�i�E����� -���ה���'���Q{��wN)�`����&�c�/�K����2�'!�kQ2{y&,8d��ԏ�F�������~+�]m�ޥ����~����~��� �Aa���	�{�Զk��:c���Q��%���(�IQ�b~�6o8CU��^��	���|	yZ�������F#Y*��]�-�r�c9�)�1_�`h�K�e���Hb�1rD�Bn�ѽ�a}=6�'A%T,j=)���X83w�d�S:c�m��GeP4K��:������� �yN�a���L���-S��8�䏔j� 菂_�+����%i�u���Q9����3<�2ͩzS�fb.���(���0p�M���!��mD�~���U���Z��G�S|�"�0���U&c ]7���(��
C�&c����͹l��R��kw��z�Ҷsw�����ώ��1�@T	^�ݬt뛘=����E�n�+s+�dZUC����JS�8<�X)'��:�>(�|��%��E:�la`L����G�����}mp@��慈 �)�5�.r��IV)��D2�  x���D��e�|������RH��tt�`�5���[�{m�����K�����Ɨ-��'y�v��Z��E��J6��,��~Yq`c�,�rI�}Z̧�B��7���BuB�7��D oh��l�]A+�%�XR�#���~N����:&���������f�ƫ��v��.3`R������7hr��P콟Q�l�ֿ<�\m����$a<����Y��θ��?���f ��fP#M��������dx��\�8�7�������!7�n5ۺ��J�(��x��Ǻ�r�]<I��Eo�d��{����c;ם�d��C�����}�شh#9Mu��ƈ��[*)=��&����R���ϋE�4A�C��iŖ|����D���Ͻ�'�$����Rʐ\A����-g��QEɼg���ψt�
���ZҨ�ح	����s	�\E��y���~�J�\X���"\��� .ٷ�AY�F�7��E;�K��ܷF���	����eo��m`#�n,kgQ� _���0�����S�O��#�C����]�.���}�R�P�Qm;�;���B�'�/*I��!<��؜�?���p���F��Q�i'}�gE�[��.C�QF���aˬs�u��H��.�GF\�6�~�Ƈ�˅'�`v\�%�����3Ǧ1E�y�;��T�E�P�S���`��� �
�d�舼S��������(���aX{a��	�I۱Ćw�q�+�Tdz�-�\�|�ev�Έ�"�m��.	��`O]��A~��o n����c䵂��w���p�ؽ0 #�{Wi=4�\-T�1����c)�I�����Q��5k~��Q@$+�HX�s��S |M5�7�S��(����G^�E��������o��0×�.��/���I��w	[��j�X>w	�d?���e�$%ʼ��N�� ��j�J?$O��CBfh�m����,Tt*�`�U_���(�V���4[^ġ�y87�5��g�J�Q��1+\�y�zB����Q�xU(�
o���ᱫmXR�7`W�=��x��wL�Ee2�!Ci�\*���#��+�eW�S/��هʅ���lw1>���ڠ}ɶ���>
�*jx�1��ӕ�����+'��GM ��Ƽ&�y �M��$�j��B9���p֜QƑѠ�*ŕ��ئy�]�V���%A���B.�a��qqy��G��֧{�	���Ii�p��xv pXB8�c��p�������.�&.J6h�e	�{�k��w��������,9��qNN܎.��0Q�ڛI�`d�~�L"SP��л�x������bs��G��u������n�5#���*e���<G���Y0�S��və�L�.3(0:�|�^�D}�����q�o��s5�K�+z� �Z��`���*Ҍ�Z@1p�1=�+��9.9�� z�p�W��&�$��µ`n�Ka�&���ݺ0̻E��@��̑G8?�}����(5�Ȗ�R�]=SN$b��{p1�f�"�\R�QdG�D�j�T$���ZJL�p�Rl����ȝ��ͣo�J���b�4��ˈ�v=;�▀�6��ŃO.�i��D�O��X� ���^g(b�F��Cx3�|;��ģ���Ǘ��P�D�ݚ���b!CN�>B~wl>��9�ô�=�I�F���f�֣��p,;�Ѯ��g���϶~�ITm~�	>�+�2����;����"ZZ�L!�[�X{v���Tq|#b�[]"�v���4K�V4�ђ_�6 �V����HҾ���D=7r�LM���,j9>���O��)�!�S�.����1�������\h�N�o��s��� ��O��!�,���S�6tD#�.��|���ߐ�"jJ�a��sK�D1+]Y.pn�����3`�RȽ�!��kp��*-@�Q)mڹ9���C&�m�2� â�H[�ZW�]�А$���4<��]%k;K����%��+�U�э��;N�k����f�+��4�W*�����۴Y֖�"��Wgn&*qW`7b�x��9ޔ8MlI�ش*@xS0�`�L�B�vӺ�7�.p8�/	���
�%����Q��P&n�7�
v�n�PL*�%�9�V:��A(�Z�r��4��(��>w� ��������],��6H���X��M��^��ؖgه�guQ3��\H.�>��zd'0y����ȍ�N�yY�Ui�O��^|IhW����w�Ѭ�o@3��gּ���U�Ŷe����G��fm�{�����n�p�@�&���v7<��&��L�7�m�4�<,�u��=�����xˎ#���RF���w�u��Ahw��V��J�9��5�5ǽ�k��X@��O��}�+���10*CR�54�zF�lŁ�T��Y,e�'��LY�[�S$˹m������/�����
��z�!^��)
���i\���Ȗ�����r8$�"$YG`���7T�*�`�v�|o9�O��'�&11���"^`��c�/�6mZ�c;S�Ւ�6ue=Ի7@���	�# �6��}�����ƀ�*�ď�'@c4L ���m�������;#�n�$�Z>�����ɇ��ǯ��D0y|���+���������6�����T�n�^���H���
�l�]���5�x:�
l+9����U��)z{$�q$����4!�hqf�8vVT�$�3�w�����
��G���� ��Υ�F��V=#fe�vdf����q��;����[z<���e��y�Q���?;B��*颓��*����J{V�fl���!�(�SZ�t���ex�<�c��A>�u�+<����jՑ&E�؆����b��?���@g�S�7�����ԭ���3@rE֧ 3<2LQ���S�����a��3m�'v�b纮�jִ�w[���9���俵E�# �rP�|�s-�Ei�1W�����`�K�9 �ȭ�kI�n�;Ql��^pj�+ȕ�,Z�%&��O�ހ��!p�O���
�@yN��m�F�����\R�=i�"n�����x��SU��Ag��n�[�O�%���;pF���Wb�J��b�=]�ڃ�>�Q��ď ��0��^�v���B�83���ׯ`�I��������!�����:����0���ay3�ԙVV�#�����u��p�!�����8&����LNּ�0�~��Ɓ�J ^H��>!��rw�D@�l�����:��x�|󐂺�Ҵ_�,?�6�4N�&�]R��r4���+
��ɤc)�j6֠+^�if����o�S���j`.��`	��Y��O��O�3U����x�UVUt���a�u���0>�~'��ac=a8�Cx��[	���R��+�m$^��$�`
�7�cbrsa�{�����1�Y� d�=���G�(U��L�z����my�qK�o�����jV�;�V�� ���B�o@��*0��Ԫ'-	; ��a7O��P�´\~��p�1�Z�f"r<���yˇ���G���JY_q��L�735$5H���f��+���B��bI�ti���Q�K���~dg[H��O��p6���覬s���#���8/�2�W�U��1��֏���3�w:��Z��W`�'��4�j\��\4 �?�\�r�>l���D^�/So�=��?���ӆ/�#;��·܀�p@�\���0����!+m�^������}0[��*>��˦m �<M���s9��~�0p����TY�U!�T���Af��`�ǝ�K+�W]!)�	6-����r�H=��$�hb�'�<�=�Q�B	#��*9K�Z���!�����曪����%�~0`���?��煾B>n�:��dΏ��Ѝ9O��$�33m{=�cϣ�[O:Ri~(����/EI�r��AT8;� �\�u�d��y�Q�;š|�fb3: <%��$۰pH#�:�@g��,�AK^΃a�f��}�r�dl����H�4>�<��?�G?o>�n~�i(�}'�]mB7:���Z��-� F�y��k��J���r���R��	Ӷ��O%ָ|&�H���>��|����",X����L�rMiG���2�݉��#��ٓx����	��;·��T��Y�r�굳�/���ɣsc
X�Q�G]e]�H�_��ZP7��`AN�s�?a=*..���I����h��%�ן[�f	-p�^�rW[�+�ue��)%S�*��Y9S	-��K�ߎ3�ڦ�H���y�<[���/��1e(~����2L�9�4�.L�ctL��J�;�ˉѵ���KL�yz���mt�v�M+����aϗu<�z=Z��xZB��� � �|� �4T��/y�L~o�����
�1��j��FU| �ۛ����>@�a�H����ź�8§b� R�T�bj�Sl�o�ɟ��~�ɮD��{N�A��\�X����C��e�F�����JZ0DJ��� z�Y+Q�1	W�'�f�4�W��ѯhP1g�Gq���F��Y�c��h�W`�\]ff	{!|�6��ļg�I��%0�r,3ʗm`A]Ðe�CG�DO��F�m����C$Q���%7�DZ�*D$k�y�~����C^ kw���M#els���c]��C�����j�A�ӓH,<�P��m��m��z��l��w�Wd���BX*�|T��Y~-ڡz'��|�	��S�)�K����������aɊ|Wi"�6��8����d^�K�&X���~_Xd���#J��t�S���\j���&��S�jI��Q��\� ��·�Z��&Lw��%y|*�k��  i���(���XUY��C��.��N�o������W7F�Bzl�3��W�˴�L҈� �?A�Kˡ���a�㎡� ���'���������BU�[�$�r ��k�e�h��z��n��Tୃ�*nM��@H7��AAGq#'%zx�E&;	����US�A�'�k]�1Ԭ��G�z���\g����!`4 nc,ZS	��R"�&����_���
5��|�B�������WK'=љ!�8t1R?�o�*�o��X��-��3Ró|�V� �59&���Ď�ÒK�r���Jw��hO*kɷ�&��M�v#�YVA�����k���*�ח�� �^�����j7�|���f���kS[h/��L�lY�6h�mk4<���`��7������:�;�Cو��(B�A�`�H�#��G���[�{���Ez��c���*L�4ڛis�y��,=�+5Tn0����r�n��B4�w1���Ćr��	W�#+SQ5���S�7`0�4���WP�z}��3UU}`#���ӥ|	B2��|��5������!�^�P	��.�AK�u�l�r̉�G��Ӽ+�?����L�?	@rw�'��=7"T�B�0�U�؝5DNԲ�=�پ�:R���Ձ�[gvI�tg�������6�D�$���O���Z7� a�R��,��X��+J��X9�^ң�&��s9YL&A�O��q$%Nb󻜚"G��Ƶ�?����$�����v��}�u��~BWQ���uH	fv�)�k�����5�$.� #ȄZF��ߛ\�I#�o>J�y➤���>Nd˰کe����]+/4�OVE���5�����pS)���\-����RAION����/R���-R<�ex���"�(f�@4xYM6�@�K�bF�-8��3L h��ڄ�F�KLhf��)mF�$-k�Vы׵��d�U��q<m��l���J&�1@o��4�  �������8˄���yWϚ۰�����������)��O�bҋ�FY�e���+�gCd��Ö�:�bO2<A.
/�{G2��0���;n2 '�w�.�U�#�Z�,u^��gT�d�;y)po�9F߽��CϾ�J$�]�uQ"�+�m�3�B%���-�[�.�� ��g*��0k�AtޙX;���&��^��>
�#o��>� br_ЯrX,�Q���^	����5�Pd���Ҋn�綦��&�5���9�y!����Uu�/���e�o樥�p��e��e�Β�9'��Eu~�p<��p���X�C��6��'=3�⬤r8P��ty	/�=%���U�e­_�D���) )l���&hYbf`�2�*��ʦ�"w����,|�_beD�k���=��<�x48�\���>�˿5�h���3j��Thp�N��/��J5���^.���h�?^91�hH�r��v�ܶ�_mن[�Ϯ������ť�QI�Zԝ	#�J�I��9� T�������	� �_#m�*��4�i��$���l��������a��+r;�~��%)�e�HY,5�m�e˭�'���t�Lo���-� @�Y�g��)zC��������*���=�.r���N1cY
)#���L����VO{�� /ۚd2�Dn4Rވ�h"G�-N�%m���~Dm,� y]���f@�SԶ��m_#���ؾY>�L����P诚��n(+0�u��s8L&��zFsJ�������h�QT�\)Y�\3[�����^(�+����{���G�įpg��}�f���xtk65b�su��,�y^�5��(�؜X�ٝ�	��Q���1<����@%�� =���EܶL�,}�=�:�F��ʲA�Ng�)�ts��V��e v�=�~�nR�)��í$�1�kZ��[�Ff8��8�!b���tf><m�/�~yF�������u��jH�N�>�<���Xl��g1Q0~�_�ȑa"��F��Ry�X�����4�K6��m.�=����23��6K��7�q�ǋ�6����e�B�x�\�S���D��)%-��&{�]�	��,��_���J���,7P�B �>f*¸\���⌼��YNL�ʉ�)I�bS�\����u&)^ :�/ǰp�)��P�d{��r�U����M�?���|Z�� M��т����Vb�Iu3�R��>ȬLghd�Ҏy��5߮P�-�|���}�3���W����I�w�qM��d}��>�:���*�rBBF!ݲ$����_9_�׍/�Ֆ^uC5�m��c�hF!�s�][��T��T�~P�3�1&)���� ���c��	"�O��p§�3 O���Z�����?��jQ�9%s@3 �8�Pyq,��ᨺ�&v�3a�M��P}Cs�C��������ST��c����I��k}U�M{�����:�],�+���U %'�����PŃ�;�>�h��t�<��?��y��mO#�5�����B{�+dr��yV��t>z��X��[��B�����������"�r�( ZTo~u�a̙(�~N����b������5QY����V�i�d�l[U\XimU���v�L{�	x�~�n����3?K����1@M���N�v��k�SB(g	���.�{��&_�Iu00�`��<�l�ϯA�|zC�gq��J��;`�4�6�(Bx͖�|���Qq�5A�׾Ƥa^Yr�����h���4:���Q����JX�Z�>��s(�R��Jf�$k}��d����\����Ŭ!L��>w�Mte�f�)�����q�g�\�[0J���߼c!�i���h����&�V��ol�:ߐ���,���+��@ߤeH�G1����+�]��n*�{���o�2X�6x� �8J��Z6��j�j�$c�K:Cy�m�U���vV=�}�;�ȑ�#M�y:;Cg�e";]�ɷK�m�+6���ц�F�`[&d#���n4I)"���5��v?���w��MlQӒz}���x#U�� �}�,��p�-0~���`=���G�v!"�W��3F��9v��l�htf(��J�'�	�Tv�D��؈�89jޜ˥��0A�`�;�p<������@���Ⱦ�=�ϧ���2K%�5�5���[EF�E߁�|���V�дw�K��ߌMm�JUe���E�J�c9U���-�ӡ�?hz���?d�^��Y���۪)P.���aǮ���9��$��3ޯz�=|� ]��F�b�������l��Li�C�J5K�L }.��=fn�ri^ǱC=^�!Tp�6�e��Ɋ�p5;��8D�G�6�|O|/������
{� a�3���� &��r+�g��:'iy�5�Q��/��CȾkr7j�e�=#l<y����AN���,�1@p^�s]ȫ����۴k��bǊ�?��>[yܾ���l�S�ϩ=06��M�pY��nO����l?�D<����9	wO�������� !� U��̑��AJ�p��4f" ��+�t�aUiaS�qlKν�p~�з/�#�ӂ���˓>���!��qⶄq#o��F���,�A��5����bl���Y0�ɟ�%�^O�q~� ��
���ϱ�2�(г�?x-9��1��ɖU} b_��W����^�S�������A�/�q�� ��O�@�%�i����g$[��� ��{�k�n�J:�ޏEH���y��C��7z��x������<g�7ý~PB�O�$�3�
��c�(T�Q�&�(�'n��5}C >Wf�=<�O���L�MF���8ɢXv2V:Nm�d�O5����'�!-닙�-�olW�^s��(*��`}��ĕ=Ğ�U�.y����yTIl!`�!+f�b�����뀟`u����=ǃ�P�l���x҃y�P-��s��=���V ��c��/ ��l$���h3Z�����*eO11�� ���(�"�ڜ.Y�Q���(,E�BoڠNwu#���q9ņ_�T4��l%h�fm���K�%~O8�^ u��BǏ�Q���`z.20�9�g����߻cG*6��퐽��R��5m�,ՆJ�S��J�5�/�#f��.�Vj�׎�����A�/zr��b��^m ą�¡�e�K��8X�"�6Ɓr-��t�#d�k�����p���T��?_X����6�s�mk����CU��%߁n�H���^uQa�d�*�V��UM��*���L��R���;v�2����_��N���\Ơ�4���L6^��a
,��3����d�E��
�%��ۼ�}��X������5�-㴅�w|�~�d�,�n
 Z��I���v�~�b4�_��Z
��J���Z���	U.N�r�-��AC�OqX�ɢ�6���Ck*.��x��������� �c	���2�m�ix �k�]��x0G%�&z��d�L�X����W�8&�����:�Og ���N4I�=�&,a�{�!'&��f�������Nڤ�Z�\���Eb�#�f��B�ӋU��C��9�O�u鬋���C�,%+���'Kq ��{0V9�7r��O&����w�g���M>��"��m��h�<��n��;ى�\��n���tX�@��턃�\Q�$	���A��"�l�yz�yn	�X �k�U�0��>��n�2T@�7�a�V�T�8���?"w[�m�,M��sAc��O�	��Jh��Ln��	ZE	`���ؖ�Yi��8�0f>���ԣѹ,��O�B���h�*�`�� ��/�� ˕I���M��T�ɛ���N����u��a*�!?y`�yy\���W\�%���U0��&�q�J��?�� �vu}�p$u�S�|���ǲ�9!�:z%& �Xm��.�������yF��*f~�G�SP�x_(ݴ����j����4��;ْ#曜����;��iS#G|�E�]�8�G��(�7�8|�����aU��g<b*�C��)[�,4ǔ�nP���!��J��1x��(T)b�5zE=W����t�@-�e����m��V������P\�k�s��6��Y�vuvy����B9������[T��5ݧ�"����Bp"���r�@X涛Q�䄬����je_�t(U�g(�usr 0���q�(xޮ˸v�>��M�]e�Xu x�K�|�Ӌj^����N�m�g6һ���v/��f���ȏ9󨨇l/�m�S����R�'T#q��ԫ	
PV��7����?S9�1�J�b����W���J�����҄F��b�M\��OBq����Gi>������LМuD��r�� ۠��lr0�`�a6"
�AO�k�H��WQ���ͺq�$��|f��nFyO9;KZS�����
�
q�o
�-����Ƹ��:���6��z����$��[޾��a_�/���P����Hkr&t��<�[j4���ʭ�'��m$)DDK�\ ��5Y7H�e�Q��C�)��	;��J�܁k�X����0?/�R�H���C�̗8|@����.��BY�b�'��#��/�R����Be��$Ǭ�ab���q�X�-Q��ɀ��SA4����R/�J���Ll
fC����L��]]J(�J5J��N|r�4��
х�U ����D���?A�4�߹৘f�"�����遉���Zr2���W՝d*��vhɒ�᧯D�������,oN����;n������+�>`��lŖ7w��NpR��'���E��
<楮���<\�2
.Oӈ��n�J�ƒ��V�.zక���%����Cv�� �@�1���u̦?�D����y�����È�l�{hZ��!�4�P�!��8�M�">����FGlwh���v/m��:��V�ۺ� ���$B�4@��p*�πdѩ�&� kmiq��{w�Ö%�r��+f�Sd�Mv��g���^k �œ�|��-��S?�I���/�}�����峘�1��֡Z\&�5
31�����b11���2���I�a�uX��n�Bt>����\wٸ�0�O�8?����� �C6-�Й}�e�
s�B�\}_~����x����XZ��x�$F��cU$o͝eZ�?�����-5�g�05�|��"+Yx������F�����Qa�	��ṔH���N�C仚J~���ۥ�Vx���&s;����~;Zc�sK S���R5@J珚��{ݜ�I`+!t�Y��Tz���!-Db�H��#ars�@�?��>ߨ$���-Փj�Nn8��d���S�!:�
X	�S��Q�K�;��>��[$]!��v���H�<�_9�w��c��Њ�(gP�Q4Yr�O�B.%IY���*�T���Sp��ӆXg�X�(< ��E]+�R�iW�C�ք�9%e�|<�~"!/#��,��|��0S�u��4�,����͙BpѵQ�;��^&r﯏�<1�6���w�p_"S���s?"�Bd�n臞G_�������~�\���!l!*��5��v,Λ�L��6r���N���Y�۲ξ7Q�Xy��n�[�&�vm�>�3W����K[,}�B�0�iY���ZG�)��Z +Mj~
0|;��<|bs9���Ð�`�(���d:_�8ܕ�Kq�AA$#�3��p������@L�_!H>��S��D���$�?��\�k&ºK𗐸���/�arݵX~N�_�L
�'G�&$�F�w���g[���g6�T<�E��]|ͦ�f�+����{G�� �=\oω 
bb���:O7�������ٯw(}�����& l��fu�K�Z�o�6]W
)�Iɪ�T +GqL	c�b=�Dq^�ngh
1�/��[�Q�g+F��틀�����0U�U��yMZZ��~F���$q�r@�Bz�N�=O�u<�u����:��!ހG�V"H?�&Mg�~oa��П�Mf� �r�G)�h���6I�VWN�vNIǙ���3���8�C�E���u���jx����e�E�Rd�o�A�w�B�~�D�<��k.ָ�g��l{v�ޟ�D��IRs �t�E�p�*)6�� ������E�xݩ2l���=ڄW@� �����秔%��ǆS���h���9h	�t$)��^D�ן�u�_qb�iX�"5Dpu�~9�W��ш����up#�G\��(塓"����P�K}�Dvn������R��8�B�V�Ǌ�f?�d�O��W1��� ?������ɲ��bb�ʩy�l��F6���!]X���:�y�;���GX����&UѲ�Rc0�f��f���&8��4\�ו��b!| n�g���خ�v��1,�l�~�Q�	��5� ��#���8��/� �l�\¶���Z8�}Pn���S-��� �7�hjͨ�N�*���=<{��!*�����l���!0�B������S�72�?�c��)�bB�2��X�;L����/�=�)V����)0p;<L�i��sj]+ZŸ�2�;0���/7G��:�M-����OР�a��b�m�T#t�qj�-����?���V�#����NX-SY�܁��&]�;N{�櫵��pl>@9���Ȼ����.��g��(Qd��9AƔqŵ�~��ML�d�Fe�'������/�Bo�((���s�q�&N,a��l7C�c�3�����%�(����/+��H����*1>��ԅ8�2�M,7om�XX���F
մGp�Q�+��'���-�R	.8��Y 	��#EcG���Sm��E#o��ƀ�D�e�kPS�D�����2���{ߒI��=�c�j�G��!����	��]�s�h�����VX��:	�Ϋ�kuzٱ����~��܉")<���ںSQ�ݯ�V��E�	��*9N0&Ň��:�{{� u�v���%׌xt�{��.9�i��2�>���:�9��}�to��6��xM@��[�T�y�xǡ��]��{�b?4�8
k�ʆ8�����ԅ�?�(�Z0w�%P�\+�P�cSM���$4�E� �d������JA�����k�J8Pa3�F�Q���՛�bey���F	_�!AE�b��wMX�r�(Q�_-�&��h6�o��n1�	WR,7��P�-1@���	l����o6Ö,��z��`��5wԏ��{��k�O��p,t��!�6%���'��XS����҉���Ls;����ʟr���B�X������q�r�M�������
�u1Ko8M�۰4Yi�m]��!�������7=��)F�7	��qI�C����vۅR��+>�����4���՝;���\��qMgg�Ʈ�<��b��\a���"��d�nr"���TLk�5�1nR_�(K�;;@��� �wV9z��c�C8o��F>г��|<�V|L7Y�C��5�>��߁;�Q�7p��*��)Eoߛ
��cߚ�p4-M��9�藾�K#K���\�6j	�����}>* �$���;q�eP
�{Vvt��N�E s�^�!2#���Q懪G��|�N�K�	���On�U�1�k&!^�1x�}��Yg~��ȋ8ǻa� � `==��鋀?��<��TÏ�[��Fmr���ӽ��t�x�h)�|B�� 3Vn-\�.��|@׋GqX �q�˱}K��]L���%��y�f?L2Ҫ:�8�����L����7��TT��\����^���e�8�w;d��� #��4�+/j�3+�O�0	����2�Q���Cբb��Z���D�/�N50�a��HNh�eʫz#A/�N��=*$���a3���(��җ�Y�����T�?-�U��PY����x�Л���C��IR?~����������1�M��U�
�\�a�/pe��e$EqU��5[`��'����u�71E_-�Y�����N,8b�&�ZbK������?�6�/1Wǭc�V��$�6����e~�eY��J`9��tJ_CZ�M���@�4g���	 򭬼2�"�e��\\ɹ�s�����,}���߆���y���uḫ�dT%;ݾ��u���g̗Rz��9�[��LF�ᨒ�Ѐ'
	�3�
�����t(0|���J,�ʼz���U�ף�������y�����R@sdC�\�˒�w>�����|p
;�sۊ�����wV���4���{k;����/�YY~�M'�Xʽ�'x�<+�W�����؍�y\M�#*0�W��EP��7G�|�L�]U�C�j=�ad�5�S�!*�}��%���g`fU�Ū�I�x�/�HZ8�������Y�y�TgS	��Ĳ�<c��8Ő�d��V�4�ѧ�K�������	�b���=�1�/cNR���@ �O��P>R�e!��}W�0x�Vy�}%���I^�u�|�"��}�{���!��|av����8<��'�]`s�+�i� �WX6�#��/�N���<�u�/37e�*�iR@��Ψ���Q��С���YjQǏ�2&]f������t�jJB%Vy��0�ړ]��iH*�g��L���F����ձ��{�oWi�TJ���P�z��w���N8P���RP�Xdy��`dqc�_읫v��zGTi�C��)�B�&a�����M�Y���XoT�xs�YsSu~�QQ�Wz?>�C�@Ѓ�kf��?t�*�T�K��|GºiP�N��0�doM�X�-ªB��"��=�Ɯ6-l�	v����P�))��>cel�4ȧ�}��eO�DFD��5��t���-8�o4�[�C�Lq��#��BL���F�|�B*�	az����ZB�m�g��_���^��
S�ɰ�ٟ�I�!�X���C���T;��M�4��r���ѷ"�4x��NR��s6��9��[alI�o�����S�v{p���dE����j��7�W��_�7P�r}���G`b�g�G�
}.�$~`S���;�w�-����ۉ�;Ɨ	��?�Ͼ��^K�t��4Y��,&>��#g�w��B�\�� g+Ϻ�����^^�6�-�Oϭl�Ⱦ��5�D�NM�7��g���^nE=��<�د��x4U �&�{�Z���U�J��y�k�I�C}�z?�H�Cs.A�~�aԲr*;v��5�º���O���.#W�ǐv�@��k�Y*724WK�Ckg��^֢�
���K_��þS�e�����,�3nR����<}������l�#����8�{3�z���U_�Gӣ	�vtn�,�$q��g��&�M��Ǝ�OYg�)���א�E	�U��B�L�;E*=�L�Wl���%)y�J���~�u�pԲ"�T"�{Z�����IZ_�R����m�V'sR%Kع{2~�H���#�9��E�b�(����4�Ô��A��/�ð�I��������6����Œg8yTDu���-*��N�R�X�R����J��Ғ��x�3�+�,�6,x��h��nd������t?ڔW�}��<�`������8���L�))D�|���؉�w��Hi�B�k�H����P"|�b��y�`�����[;�_�������9�t�h*Ns�Mh~�9�+rn�v�5�)�ry��G}==m�����r;��!O�K�p͑ˣ�&0��� ����j�h�*$�b�&s]Ԅq�x7f�@.D\bCRylaF�I�)�N0�Ч����Q�.O�SIZ�\a;���\�΁��j,��J1?��{� R�0gA��kvƤL-	�Rj���8��p�poc� \&9��Ðx��[��~�Ţ����U�T��
���)������i�f<x�|�IbGk�g�]֟V����X�m��՜�r{iFҹ_g����*suõ�-�� �o'�U�,���L'����.}E.n*cC���$s0�/��Cn���*�W�q���&��:)$���_��Q[{C��iT&�o�x
3��<�9}��ǲ�Պ�_��#�����m@V����UO�c55K��خ��4OZ׆�Si�h�g�y݇ �z�̡c\�5Y�T0=՟j��J��ϔ��:b �mM���s�a֪�Y1hS�h��oX�z�������U* ��'1[w��PhhPyI��n�-�)�qk'K�V�1]��	��l���#��"8���~)9���f ;G<0�������!Ë��L�B�I� ���&�#�ԁS(�����r�k
K)!g=7�x���?`|)�йH�6�p7��w�<0��`��B��g�%�w�̊ 	�t�.� 9�S}��E:]����j�����S��rkT���˃he�w�B�R���zuh͔����l����D�ͺLb�R�����h���J����8s������cg�.�i-`�µ��P��V��QЯ%�E���6ɚ,�-���.<aY�xS%_��淪#_���H<+�����ʧ��)q�~�����`�>�;s�鉧F����5E��م���W��y�C�1�C�������W� ;01V�鸟�~\�Ϲ.tVj^]u 8Y]�XD�=T���H))��5<f��OH�+�w.t�|AO}6��x%�3�
-j���+�<Cժ~Iz��˝���νk瑦��oY��)��L��cҚ	���Qze☛de��E�Z�d�M]�V&��n�\����\�^���D« {����j�����a�F�BLb\�tK�r��&��r*f����B���+���^�.�bmis��s�C�C�b��b��O"ͫ	Ӡ����0��^�W�n0ϓ�j����B���c��HE���/G�L�%Ԫ�.�=wH�_��u}zz�'$󡮔 �o`�k�7��ar.�P���B��P�����p)T �d���͖�.ʯ�݁$�2�6N��R��U�r\h���M<m܀[���z
�-�Vd?=��>����P���]Lpw�a���x���˳�h����.
���k�ᆙB%��k���Vׇ7����9�;�<]3�<$�]�����Vr������2���y��>�0	N���GJQ�ջ�V�����?/S��L�.Rݨ.�Q7S�hj�:�X�{U��L��IT�>���E�_����b�Q2:Yu��1����N;��g`%
���駮��,���dOd�J+1r&T���}Tj����P���JʳOwl�.j�S"�Mz���x�*�'q_\O��J�Th�քk�U�c2���|��Ac�yڎb �����������*��ֵ��T�a���8z�}�!�*7�u�ٴdoLP��zA!S� k�覈'��9(ȡ����y��H��h�<��/'Nx�:�e��K:jWH�ψ��ϗ'�X�qHv�M�53�7�@��nȑ�qϨ`�N��~ӆ���ձ;�W��U����E�c!ӁN�-���u�^@�x�=<܁4�E�d�/�YP�I��S�׎�W��Vi=|>�Nr\�mV%�� h�G_)���~��b߭���"��&��{]��\�'0ػ�{N"'���$�i΋�qY�?z�Ѵ}����V�}�R�n�;0���Zh��w�޾qURwZbBS�mt����aւ��ԮJ���as&�(��(S�Եn���L�v>ZZ�Q��"�N80e��w���k�Ϲ��?���!`셽4��b���E����O�<����,휴���I�2�ت�L!ȫӄč=�p��(�½QyjC������H�^���l2��߭(o޾:.+�Ѷ`kW�����Ɨ����z'ܯ�Bנ�dL�U/ o}��)Ҡ�~Pv�"�#f [V��"���46�%gZ�c�gm��e޷��;HRߠ�
O} ���@�=}`�GK���)�Ŋ�m����v_2����- a�'���P^���
�����I�(�'P1�/6�P���w)҅��L?Qb����s�n?��9��pҴ�����+EW��76p�� ��Vd�\��5��\|��7A]/6C�Z��7`x��)(��H�ǌn!o�}*��Z���7
���%��~�|�8[j#�yM驓y%��TwGw���	%��Z��z��Z�oLJ1�#��J���:%q�O��Rx6bEq��vHAX>�+UT�"�1��ի�׃�v^=ۅN�Eč����͓Z@���ȃJV���S�Ɂ19{��-�:�x��5�=��h�@KT���դ���`�
��Q�E��s�"�c��59�t�C��e`����u_Nq鷬V��m�������jH�I��_�x��)o'ٵS.W�2����7��4f\Bo�j�l���k���-K�����XB$
�o$��,~"|�y>a�т]��LH�FR��(Z�JW#�Ԯ����p�~0��P6R�Ul;g;�DS�e���mG�A.};��r�ǼǠ��q�(��$c�QH\hJEp�t������XB����|�7���9�V(ַ��؀'���]J��)c>Z��C,	���B�f:�ݒH��:�Q#l��Uw�b��%k\�((�k�����_-��	C=����뉤�:'r���Z����u|�:�Ò�|xJ��ļ�A�e�fU,��J��H��j�����A��`����g�׈��^AxX��A�Գr�� Ｃ��:��6��������#⯽�N��]u���R�������s�2aU4.�5��YE��	2 )������'�7�$!��%����q3n������mjGHɝ{7�?Aq��	ް�	���|���	�E�=���׉�d&��R
���6hӟ��[>J�_������W�{Z1��w\�K��oɖ/��|����i@kc�9���=�˿�ȩ�7C9��A�L�Q^,�d�Hg����έ~��Y�����BU����V6V�Ҧ��--6B��%	|��Y��*Mh��#�3E^H���c	v�)�l
���v���;��߂<��D��h?n��V;��SHw��lѓ�F��2�	��ծ_���r�XiK��[���1����o=���š�6�HyE����1L��q�����n{m�dޞ�X��5�FN >=���C�rg��v�(�I�N7��pl����C|J�I��n�p��,f皼H�X)�0�J��ы�I�ކP��5>�0U�dg�bs��;����C����HE�8�;�E�X�ù\Q��tW�楪=��C�t����	APX{���>�L����UO��Iخ.Z㘟q$A���K�"� g@ەw��^��:y{6»FX���q��׬	�Z/r���t�P��ܤU��u���J=Q�<8T�v�L=��O�b��s���$<;�ѩ��M5(x�!���	���}i.� C�����`EZM6^��,�?�~$��Fզ��ϒJ�2+g����u���>��w���H=J��;^yة���+p����&����ɉ��T�g�T!
i0{s�(8�怉�$��"�O.8xf"Mҋ�s�?�@����\4�7n	^�L���>'�����i��}cQ�e��Fp���ؑ�m=�[���.�����ۢ�_����4}Ϳ�? U,� ��,�c4A�~�bݛ��%X���N�mu_��3�u]p$v{�~��z�4� ��X]mך	A�p� F6���:�s��DH�G�Ӂ�	M�*�R���|����W��w���
T�O�DY "�A��ڬw6�I�F�X�$�5�q�Ř떀x����}$ �7j�� B�W��������?�{b����(��ս���Ie��(#8���1�h���襷A!d��q�dj���ϓX=l����{��������$��r��>�K.{�EJ���Ƞ�m�~G(7��Q��C��{�8zl�X�W3k+��"������å�M��n�g��U�H�S��2���t#��Ϛ����[�E�9�)� @Oa�pp)=`�&w�bX�,#h%�S&?���,�F�J��~?�}.zO3Qxlp������o�o�dc��M3*��YZ�^����h���I��a֯U��ܱ�rr0s�rUgMkʷl6`��~�ы�Z$��dl�d�J���@ƞ*�5�6]��
a�E��g���lp�XB���;�F�3Ss��;r�*��bPy�j�:�N3cDԿ;�K�x1���$�:��n���c�f`�0
KG���C��J����\_F�i�Rw{���3��g��)��Þ?U���>P��m�l�H�d��� D��H��������Ə� �,R.
�ML��<{;s�	���G\#>�����+=&�֤�V��. ����
؅b7�$���a�Ω�%֞�a3� Ơq���<�i��з����	~�)����N0�}Af��x���Q`�r
��U�Tt[�B�JZ��L"�'O	;�0d�H�~������\�
�3�ֵmS(�)�)NЮ�o{��U@���ž�\�xK����S���76|��g���p�O.�#(��<�,�-���o>�~���Ecuz�|D��>'���/��Uص^+B��GWo�#���s�G�+��4f'\M}�X�)'V���}��ӮrB �/�$�7�;��2k�n	��v\�av�.|a/��a�<��J���|6)@�3�!�������z��wu��O���>H���ʫ{�N���6�"I�,�i�
��{Ǵ i�M�Z����I�5Ӆ٘���ĩ^�&��w�j��&xǢ�CZ }v���Y.�l$�d�kZ��E���(�ߘ=`�w��?�Hݕ<W���5��^>g?c��e�iT��f��t-�ɼp��W�{Is��������:?Jo�xu�aB;�x��M�;N���e8�:,#C�����RD]�!�2� �G���Z��5�t�Q�+�Va�qvi���[�#)���^�����{
W#5L`����3��2�����ҽòⲜ�~�7T�XJ��
<��4�g�f�m��I�W��$��Н�o�� ��^��ig1��kJd�e�|�޸)�����s�	���_W4��L�@�U�fQ˳m�V�(W�K��H��L�!����%�+����2)�d1o��fhK{�XRF�}�����j������ѕ�����J�����0TZU��-��QR8�Dʯ��9�������q�fT�-ҵ&ʖ��ߓ�O"rm�z�km���g��;D����aր�m'&�b���<�f�(�6(2&}����-�m��q��şq,�g�9�*��ʵ�������"1:�������>95jKH?��3B����5���{j8%aL���i���JdZ��Ɇd���N���&�9�əD�WM;,�l�n����Qs�3M�#ߦ�
�+htH౳��BCH;l��ׯ9��X�?�C��jOz�G#˟)���&�PZ��c����a$h�wA�xh��V�)��L_<�s��,�F.8f��kH�gk���B�Z�GZj�r\� ����D�A��{��/T8k�unٷ)]���o4�7��\8H��M�|��C]�>�̃d"Xc=�����r}�������7�?�8��9�[Ǳ��!1�]a�u���9k?`§�����Z�j`�N��*��5�pKY{C�����]�B��V�|j>Q�����(�X{�� �b�t$��׎j=*^�E�{Tp>��c9����PV8�9?F��N/9�)�Zkz�s;��')W���A�vǹ�4W?�o�u�L�!TPJ�h��8��6�_D�g�]^qGK:^��<�_��[J|&�qDK�Ď�.UCY ��zrs&7��HVܧA�Se��q��� ��x�b*���6�@aX�|��� �������ݜz4ΑxY��2��;����N����l��*B�C�[�c�8og����©��/λi�9��d��#"p�U�GS�&������U�_��؏���2�r��Y�6�q�a�688S�ū~��:�+�.�Is���������S�̑
pz@?�q���P�^�/�l���7m�����{&7fO˵7v�i�d�u����%Mx{�Ҡ�;�Q3�y��}J^P*[mTӰR��5I��wL��}'���Us���v_���2�Z�HMl��>B�`���(b+\������~^���^��Y��$��j����;�[z��ٙ�݋���W���q�J�77H�!���'�M�K���Tn#�a)r��l��l��	;�%�>$� ;�ŗ�i�O��U�KQ�J������s��mǁJ.�?�d�zP���h#��ehC�$\,��ܖ̏!��/�%�Vv��1#��x�UT�E��%���V��5���~f�w��b����a�p�Ҝ�oZ#��p��fB	�%R�3%�u���k #�l�`2/�z���Y�:ۥ�Cg���L��$.^�򅤰�7poH��Xv��\�'�l�U|��C�{8rm�!|�tN��:��#����K�� gw�a̍4Y�9I�����(��z)�T���>�D%�-��6*ȍ��R���,���X0��h6ґ��v�`��d�)s�m��;$��z���ۀ14��I$�?��������MH���w�����Y���=
�Sm#G6�vW�! e?�͊���k@X|G�uO�g9+�&�4!�?h��w��.�p2��t���X�[�Sá��4-�@�P�Uu)7~���@�!�F/k���X�ꁋ��W���<Y5\эx�y��`Ð �d���3��W, ��#lɔ���I��Hk��j̣��3�t�]1�r�]���>��W�ٻn���N��n�wWc���'[tQ�CT�>����{jU	�谰���;��ظ������KB��'��؝iR�!�8��pF����0���U�{��>I���є_����v��[fk-�gtf��X�#l�"Y�ђG�@b;W�g�'F�aҐ֝��ڨ�β�H�����?6�Do��m(ގ���d�����R&�1��#+N?��46�ȥ���&Q~�� �d�N�Y�jdJ���$p+7a� �PlO[6��'��"<�Cm�bs�h�O6�d�ٲG%���-zL����ЀV�0XVG ;
�vA�!�
�L*`]�Lk=/H8���7��7a)�U�	+�mƽ���AW�L����P���8b�Eȑ�K�����gՋ���L]]ݥ`���N#Σ�8�����*ZZ<�sM��Cz�jo�nip�{�4#�O�=�[���<�z���A!ճ~E]�
�HQq1�%�~���I�{y�T�p�+����K"s���9�����Ē��%���m^�EP�6/h9�9��3z�
�\1:�h|`�����X�`UF���3{���Ad<��Q��z�4��~�~Jաt7u�u�Dr�
X��˗��C>1��dAX�y���Y��]��y#o���$���Oh�nG�����,?�vI7'V~S�U�&�2?y�

���i7K�@�R'�ۅ��S7��諟q]��
m��$s�x$�}C��V0
l��EͮB��j�ڍ�,�2�NL.�����6�rXP���1���s�	K���y�ye���v�;dEj�|pp�\rh����\Ve�8S~^�����t���+]�:^طi�l�.��1�]�.2s�r�[�=��5kL��%����C�oCR�p�Q}^�[T1��3�&gC�C���4�~S>��*/��a�g"R���`y=с9Z�����7��ԟ�]gnM�F�)�Vק��𨐛�M�~�2����9�*;b
�^ԣ��4~������D�ht=7����}lB�����k?�֬et?���2��uІojS'��@�
�KP�E��
Z�t����8��L�1�I��a\p6�6#�ݕ���g�_1�2_�����A��!��������'pϯ���"h��R�gL��e��b�XTp��$r��Iegʏ����ġQ�����u� P=#�{���8=VW��V)�s	��4Ʒ��˵͵��r�gnd�bt���L�Y��i0o2y���
_�_@'���p��y5�FJ��!�������Bl�����h�x���L=F�;�꫏�D���w��KY  U>8���hx�����E4$dϜy���-����"�T����qn �e"�m��`�,c�Q;^�5��>_�u������1N��`��rlD���h__?D8����` C�����Q$��eP�YC8ѩ�U�&l��u���
ګ���8N�����P^�݅Y¡^���&�&�>�{Bf�>W��F<g�2C�T.E��и�,pj��lR�v�YPr��;��Ѐ��[	�����Yר���[�<c����3��{��+܅���?[��%2�a��lX�ڜ�y��J���~�>\Bކ�Jy���I�6�~�r����R�w+�������"�
�
��n�&}�5&0e�K�w]u���D�ѧ�i΍ݕ��O)vѣ���B�em� DU���N�y�s�:^-=U�*G�#�Ʉ9 ׳u׌K����pK8��V�H6��A13���ij�*�?�������j3�����Ζ5�ѡ�pGI�����/r`��_�?�0ߌh쭵�O���s��ŨY8F�~��)�;��F�����	�PE �O)�}%��y6�3	5���n����O��R�(��G�z��ɗ<�j�����gp�51!��c��D]�Ē7WI�������Z ��^�"Yg���C�	��7w.��X�^e�^k�C,٦rС%ʲr�Ȳr5�'�a�i{�"���䒨��N�4H��%��'��p	H�,r6J���O=?�Hv��
jk݁I'�nY�Zn�n>��/'�6Qa)�H�M
3�_�)��AU��������
8cZ�m��}H�N6��!X�f,#,ǣ�-L���`���?Hd�iK�
�d���S��(ܙ/����Z.�|�H�g�:/��rO��+i'[<��c��n����j�Z�ȥE��1*�#0֕`�(i�?�-vQc�v&��x����H"n&0|���T3��!�����f 𐋂�J��,�E�-���I���#�#և�£Ǣ�*��a��W���ʕ��Ha�¦�E?�����BR#�] �(F)j�j��S���q+�1;zM®HB0�ц�@����8�����DX��2�U�pRF'��4�r�wU1˛-:Q��m�0>���s����%�o$�oʵ+���u��qV[��� �v��a�(T��_�z�E��fPC\	1;a��{�A�Ƀ;s��p8���ȶ�UZ�[�2a�D �!퓆��-��%v�![�:����hQe�Y8��7n|��W;ŏ��a̖]���0w��f��NQ;ʭ�:%�]}�@v���C95�|f�`xĆ�c���˲egd�fۇ�[*���QM�Z�بj�t�F5�W4mAR�R_�����)�/I�FXC��[�&��}-�������1�����(->kP�"�'���qm�q���.�l���Ո�*u��չ��9�J�k��x;�o�0�媻�Tȴ�V�z�[�����~�u-D�h��U]�?�Mδ6�9��Z��D�ݖp���'�3�F��yK�DSPɞ�9��U�����sf�ãa�W|\Ȇa��D#d4�/k+ߩ��K��#O����HO�ִ]!X��5�]��w������A]�!D����^=4$�S�QD<�l����
�u׼l� ����߱*8U��l5��9n���c�,�m8����ʕ捞%����itԟȧ\�o�R~`�֓���p���0{���y>}K�Q���9�ҬU紼��d'�.>"GN�(Jgr�����ZG+��G�n@�cv(�04��]T�N�R���Ā�!�.�2��cc�:��0�E�k�+����2=%�����,h1�	�эŪ��+�6�@�#�ب+EM+�˼0��Ի��m�QS�Z��ǆ���$�!���D���6�a���$�G�|EIH�Q�zj���j�,w���i��h���Z���i^�{	�ekvM
G�F��E5F)\mK-;w1����؀f�x�|��]]�V9;�)_y�G=g�\8Y�K����D3�)��=� ߄�J�K�{NN�Qj2� ����g���a`O@qt�sD� �m=M�S�(o��'&�t�X����� �@�,&t[E��ȯE}�j��*�?��6��m�躘��0Y�c���ct�g�Z(�`��Rz6�rJU���T�"m�G���SjY����@����=� �t��h�>~F~IҞ�b,���4�����$z�ܹ���s��l�ܢV�	;W�[@�x�6͘�1�g��=�ڳ&��a�?��羘G'���M"%�}PU�<b�<T�n��om]������k���r�K~p�WH��Φ.�RI\��Q{_1k��s=����Թ�ΩhR�J;U�EYq3�~��Pw����P�nD�.GP>�F��K=e/-ǰ<j7��va�"��.�2�D�.�)U��Afu����7q��/�f0"\��wiO�
�	�������h|���2������m�h���g:�^���a>�_�LCꖤ]�
�<��\�^7��ex
��1gEM�����z�+��*����ɤ=mM+���׊�Vn��ϛ�o[Z���>i �mb��XCOoF�;?Q��=�1dI�YO�H�O���5w�!�0m`�t@���ךw^Xհ�v�ۯ��Va���9Z���~vxLBޫ���Vj��ή��-S{Fu���%����oum�m4���CNn��D�s}'�s��lh������B�����T�ꍗ�_��7�.FK�v�XXu" a1�0�C��u���no�Mf�vK���G�6��m����7,n(U����d���)R�Q���y�����S�p�+U��ᛦ��&�����xW6i�оwA�.��4T3�������/���o���s ��h;>��R@�P��{Ǒ�RU�}�}e�ù�c�����j��3�J�m�&�_u"���݌]�}��(�H�3cl@��0C��A�O��0Pz@�;C�XI"s{��w<��u5Њ��p��iD���>t\f��K�6��r�5�	6(If)�lesU��Ҏm�3�K��x~fE+Y)m��hF>�U�8�� s�@�<����d�vP������G��G����^��؈�9e*��:3���t
��%���dǇ��WLl�;<k>�6ܸ�CI'�{���r�,;��D�H^������(嫠���j�f5�d��YzH��x��
C�U-n���[#o�u���ױxg��}�eU���Zae2rA1o�]U��N��O�تԫ�s�l�(���n7s��B�H���.#��/C��S���mRE�"EY�4�����B���DZ��f�'�Y���"�PI�;g'dO����`ͳh�@_J��du+�8ŏ��/\T�Q�1n_O�)�spC����7vd�O0��;�{���j���A[�"1M�O��������_
�mF������,g*'��JE�eF'����!��y�җ�����d�,f%�UC;\Z��~Z�.h0 ��yc��bp�����4u�e2 �H�06PTVRNj�(t��Tg�N�pO�[L�+Y3���5���p�6�48�:QA�n�oE�.�9ʟ�g��ꯍ7������i햣kG/�@e�M��a=���{6� Z�A\<�� '�h��&/1��5�Zw�%(Ԯ��0մ���f�l�ƈ�1��]a̷��A��C���
h�c;��ֹS-h�4O ��(՚SBT�0Z�%���R����<��KoF*8[������E�PC�f�T�&{����Ur���Ғ8Zە�P��޿�μ5��݅����L�B���[D@�")�|�ڥ��EK+�a���<�1iG1�קo_`�ع�=SwJ�z����0a-�'��p&)	녀 �������@V�Fyq�(����{��^�-�eᲄ���m����x: ��bb�f��|�6%�� �
�F\�,���u�X?f��xn����=��Yh%��X\ܰ7us��ytX���90k^ x Y3��v.�:s�Up�~�m��y�ԌY�$�8��2���5�Q�i�;2�@��n����7f�G�9uE��X��tv&�����7��/�2O�bIPvb��\�B�sV�C+?O��J<��w�%9Yz᠉�������l�@v�yV���x�rh���I�ٌ>uJ����7���OMeI,.W��X]�y<"�����W�������G��S���'@����k��?�tܯ{�7��oXq��4,�B)s��6���
���\�,�M��$ST����J5���,m��4$�&�n����e�����|$��ϗx�q-��8#zT�\`���J�2M�1f/:0�mY��L�c2�Q6w��>���F��ƛh�����:��U�亠�*,�jNx�T{h#Lx+�`$*�V����ţ|`u�jVn�!l�КV�9�����(��!7� 6:�ې��\�_~�f�(O��~_�%�HT��m�J��rt%�R�(�J��k*��Dmm}:2�(��ߖ)X���Aޝ\����,n�&���i.�-;�~��X�6{؉
�s0 Q�Q=��	8ǚ��P����g',h&��������� ���ɕAuV��N�˘^7����GE��SD }��%���v�W�01��f-O��kv�;����Ӧ
hʽp"���x�Tq� �'��5kr���,�p��1
����'!WvtK�0$*8r�꽀��%�7�T�6�E�,����U�h��$���d�H�'��Ij��"�qH���3�\3e�ۗ�æ�#/[��}�	��F�E_���o���@���0k��<�U���w��+j�n~,�	�\���4�n��a�p3C6�1��԰'������x+o���u*j��e\�K�b�����1����n;
��"XY�
�'^L���W7+�X�.�e<�S ��a@r�s^�����oL�:��2�����'���?�*�%]a��ѭ��=�0N(���qYo��N��g����9��b�/�.�=�|��,����I3m��"��d�Q�_�g�l���r|b��a�M͠T�H�R�z�t�Mv9��|��lqlCr��u�!t�Z�t$�p�!9=x�p7��.�z2��dƯ�C��-��KQ���f}�z��N$t\Q}�����y=ޭtF3{�˹��&�盉��� 	�hxw|Tًf��+f���/�O\t�s�ȟ��=�����r�:q�tq8��� 8�I��Rn�<'{�A�L9α=(G�F�<P��n����? wc�r�`�*�;<��{y����č�,=?����"��{	�/|?��<�CT�4r��p�q��G2�1}����ə�ٸ�������I��KA���YA�7������|^�����Iݴ� ��T���j|�3Y㎦0���qTB?�G���N�RQD)B�wѳ`��!��p���24z���\�~��{	��s��d�.�1W�l�?����5�Qh�Ν���[�k4S?�l$��eI��q����aB��C.�?�[��088d��dt���4��#���8��e�ݖ�N��2���	2iS'�@�J�Aj�\r�t�z�|��Ґ��$\��m���!�>��Ig,��,/P7R�D{'I���B����\�,]���٣��gBEQ�4� ������he;�G��vO�[��x AQ㋔H�w2v!⋏g��X���
��5������(�0���3�#*G�~�qv�](���ӵ�e�kNѾ�m\��
f��+�]l�NՀT�Ab+��M�I�q3������ �q���I���J̑�͹�;�u9)Yj�(4�?���a'�v�������I���!]Qۜ���C�6�?[�j�ɺ�)�J��T&ЛCv����l��e�`Nwh�f����|�����l�1ޔYܨJ7�zt&��Ƶ���1�N+�ʵ������T*��U�;٬^$:���$ڲ	��^����j�5���r*�\}�
�߭���M�u�^>��òh��s�)xF�7���^Us����6��hz��2�*�M�h!�p�L����:l_F�w��~�V�:�d����e�@Q�d$H�����~�F��N-����$�zDb�b;"��@%4�򦦫:6t�S)ư���e˴窤�ƿ�[��	���PDk��Stѳ��H���,W�S�4sJ�d��\�UK���=�+,��P%e�Eh.�;��`_���%�f.�����̌0���  vȩ��L���)�)������rI����S1��+5BR8�ל�L���F�Z�R/vh���d�R$����~����w�@H��D��<ZCf2�r�R�P�e5}?Ѷ��yǗ��`���Ɲ�&��xf�+7}�b^�7������cu��i&_V��8˖��R
�ǧ�Ԥ�L�����	�$M��D+��-�7��g��r0Lo7{��`~0!�W�ٯ�[\L�2�:�"ڻ
���y�Y
>���@lɪ��@��a����_�<>�� ��&�7'��´#���o5܂h��ц����<�g��c���V"N�S�9 ���d0L�Ӆ5ȿXlY#��f�D�����̂z�Y��P�Q�Z�cg��K!K�X��}C&p6����F^�Ã����`� �Ր�?&[o��Ӧ��1�㨐		\tQ:��,��->��̘j8�$ZU�cX��J�Y����(h%+4���
ʵABx�_�&�u60c�8|U��y�8+kX_��6��T���Lr\�Z����u�j�$�ϼH���X���&��`�6�R�1�Gx��C�d�L�ͨp����F5���h�v�"{�B!)�q�9�o�����w�+���	�m����}�����;�\��\OVc�L �u�ޝ�c|���؛�d�r��E���)��Hs��krl{�]�~��c�siGѭ���N�B��m�d3���"wv�?������D��l��-�B�d�<�� ���y��dfN4{��t%& �W��� m��A��&7�0,���7���H/����dZ�	�Se^`��$a�#�o�Z�}�lg����'�����w�ڰ�E�O��p�7Ӿ��ͷ�(T��T�����g"�/:ុ���/l,Z>�=�����7�v��E�A�t�&���;{��6���$/R�W�e:uA
��x�������+T�S�4]r�#�>�̶��g@��J���ϸF���TeL8ѩ� !5�fƉc
'���(��P��?�n�1�d+J����;�����
�ҏ:C�.Z6	�WŚ=�%9Y�o�xk�.�F&lO?��ో�d��ϿO�i�"[]T4�1P'�|ʱ��h�G�=��Ĩ�`�Phh��S�Ƚ�C2��������x�LL+�N�`�~���j�F���g&�E�����
��
h\�F��#�S V8z�&���{��S����7���s(+���]�i@�wt�TR�<%D
%��8�q}>\E�V���f�Bʩ��}B�^#Vg{���;@�ܔXes��~@ٍ�&���� ��'����U��2u䫏ܼD��#Hw9���;�1�G�T�M�з]���'_ᗎ���\�ˇ��y�n��\
��S�j:�a�caD����� 7���.ib�L͎�@�j�9��HlT,!(i�x<�Wq��1�&��Q�� �]���b��p� ~�p=���I�5�+���>�z���t���#Tx���'��,�A2u�3UG?ɾ0�3�H�?oQݾ��0�j2hQO��]s��AXr�G�ʄH�஧�m�Z-Q�"�KB�k/-~1�p�4\�/j�>��]���mtgEB^f�ᒋ�\N	����{���$5�����T��UKy�.�a0˰�O�/;�5[o��JaZ��Җמ�˜1���sV��Ʉkdf7����ti�����(b�Д"��S�LCވ��/�?��E_��S��B��K]����=
-9
�|����Tѝb{>�^��H|�C��L�-ֿ�.�Ǭ����gU�]u�1!�FDvHyKU�����_W,.�� &]C7{�|�����;��u#��lXt�����R~عX�ן�f*'A����^ �P�ɨ�<@�v�9��4S{�Hhg�G� ��ܔF�����������''4�O+��&u蟨C#b�b�L����[���?ݩxE/3n"���`rH�ޏjY{����)说����o�g�g&��4��y����h����@����д�?��c'�.�|3��X�z�(���F$��f��vʼ�fz�9W��VC)A���AH�L�M���`�n�4��2+#^)
x���Pm�lV��L�NX��'��+��a��)r,�T
E-�ψ��w����E-�ʓ�x��h]�e�y��,�X��Yi�7�q��}����qfR�Ω
U.Jn�e���֘mE��!ljPB7�~�	n���9�¯�T�$�G#��Kf�cji�ۊ�x���C'�&P�n�כ�Ky@�i�T��Ǯ�T�;�>�g�r����kT� �96�*F_����w���J��	%��y��|�pO��%���z i�h���$���� Zv4u�N.�A�EDMqZ9�H��6Y��ϳ��_W�ߏ?BL��('�U��}���I:A$�IօDr#!6V�k�o�� ����F���asŢX9��0)�>����KY�X��:<hr�U�1T���x������F���o�c�n?6�CCu�4�V��:W�<`LL��x�
��lw���Ȋ[�)	�ڵkE 3��%�FI{^�ul��<7B��g���g�!n�-�5'�0���b�A��q�I���u,C�����*�ϱމL�����xO�hsNB+�XN.�(�,�W^������\���0����������愥fp�x�NŢ	��i���1�8�W0A��\�4�2Ǎ�5Ѧ�#��z,�%�O��QK�օDЧeQ}wvq�u��iR��ڈ����q��z��{��t-���/7d��![���e<����0}� M�܊���>��X���"���9��®\
�.���_����+���샍\��X�\���$w^)}��a7�[��� ��0,�u�����1����C�;�'瀂.�+�,�t߄c ��M#,�C�ࡢ�e^�^K��S*㭊In��ς��Z�K�:o�H�Ve�l��#��Dnf���!6�s�� 6�c
���&#N�)hZ��T��`6$��Pt�!DF�[�����4?!b�ܳ���`MB��e~Z[X�D�ez��T���q���~�.�B��[�B�N���&w��d��
�/�.�o���|�n� ,a�$�:���@��an�G��_W����ɝEe93g9�!��ㅣv&,��F�nm�$`�#8 ���6��I�Al^
&2p���:���<C��.PA2e�w���}/F�Ƿ�[�-�ߣ5��� T'��I�N�.+6n~$$� � {t.��N:�R+��vٽ�f;.t;��e�B1�c.�SIP`�(�]o?ԁ����=���s�?�����5��;[�H�)��F_zl��K$X�AM�m`��oz|��:�Ohf{�╡��
��*T�T*D������L"��H�\e�}o�L�;;���"��g�c��T��J@��{����5 [#*�r���P�S��.�/���[C�c�܊$$�·�Դ�e�\��GD#�
��y��)�(l�P*ƃBU~q�&��~���J�ϛ�87I�[���z3E�Β��M(�ʣ�}'�Mo),�o�u��
��V�2��w���=a���a��q�7�_���I�����j'��B�iz�P	0�$�'Y���|���
��9��as����|����vƺ�����Q��/�#$�5Iy��5N2ɥ������)�_Iq�1M���M�2�z��)(��Ӣ5���9\��b�5X��}�|��nKA�����d�R�1\�2��G2��tS%W����B��؍���>�����w�*����(2}Z�A1J�bm9p�������)!+����YT�|��B�zFʸ��y�q�p��|��&y.(c5ǚ�A	A�z��n��/@H�}�<8_�ay�^�h�G]��k�(u�0�"��b	|�lS�C�Pw���$�7��vÿG��L�@*	�ېMyZb�R~��{N�i��������G����٠�#����s'�=��itt��K*��vT�
M*b�2eD�����'��恢��~:Z2f����V�]�@$�U�R{gQ�8��f
�joX@]v�'��U֕r��xڡ�k+p��w�+�>����k������>�R�uկ�,�Yi\~_U�}��.��}z������H���p�u�>����mt���y �%��̓���/
a�>mRbu�����O������nU�����#��l Y]��'^���k���p̀J7�0��nO�~�p�\���Y����,!Z�I�g��i\��^1�*Y��3��m�t�B��X��d"i�Ӎ��kDCp'�c�HKb����6����|�8o� q	�d�>��xRs#4��|e�ę^�h��'}�Kb�=�&�q�ڏ�`�9F$��~��v���ޢ���=�������0^�b�t�����H�H�^k�ݰ���(��ӛhK9��NR�9PA�L�Gq�S=C����s@���'���r�T�k�#�?�]n�����J��8O4c���g���}d��$J'N�u���߸��ӿZ�(E쵋�x.[Y��<2�?�K)�並`C�ѳ��S�M3ŝ���nJ0@��'�wB�����Fy�<��tRN�c�������0w�?(�њ��٣���:�`56�G)��W#w��?Z���&�+u1��"L�8�
����-��E�*�V�;�YMՌC�M�}�<"��+̦P�Sh��6�'we-L��nT��&�6��[�ȡ}j���iΓ�hl%��V`�u�ᕄ5@��_��pFʽ
���1P��8z�9�Մ����p�X2��ח[3�L��tpW�k�Dh��\���fۛ2+V�53���7�?~��q�נ9¸��]V�nxU�!�$˗�����D5L�1�*+�h4/��[/��Y+KE��hN�2�� %t�3D[5�ɭֽrr�1ǽE�.�D��~}���Ǵ��}����Y��`��,�)0�����K,N����u�/vo��`�i����
'"|b�Y�y6e�%-��Б"���c,i�@'4������/��5�Xu��~�Tԇ��kȂ�>��&!F��B �X����1��*��= F��ޜyV��k�g�`��Yw8g���<�[�\2J	s˂Z�\�g���VP2�)��s2h�9�����:��or$����5 _�`<aK� N������2�3�6H4u���sN�Ɍk���B�Z>/|���fbW?ѫ���wV%�sx�I�i}�h��v�L?cs�%� a1�0�tx�r�Y���V���y�\)V�]r.�gt��t̙�} #ĕ��bl���݁C�{JY�v�t#bF��)qk&������a!�Y�*�K�yb��A!���8�O�V�(���?��Du�����Ik��Wq@�׋�%��P%��@нw��Ǡf�*M��ΗP�2V9׻Q-	��Z7�����3���|p\#��6��x�>U�_�;u��)�B}����-vYD��C���&�-�~T�Hsn	��j��,�<�x���o+c����<*�h|C#��
��7d/�Ĥ2��)��F����V�#���gt.�R�$jx�ݴn ����,���"���<(7,�<�&d�ɟe��.h��
�V7˂��3ND���L�9����^�^���m�X�_m�rw�����<�D`�)8�靾��l�d\������<�H��J
mJ?������/�+��Kh+	P�&5Z�:}<�鶎�>#��Cn�YA0���Wc��6)�!t1e������a�'#�q/*� .�ch MV|OK�W1\�Mp���YJ�h�n1�"���,B�`�P��4� �w5VǸ�ff��Y�QXL�c�o�6�	��������c�����3�����(��&�C�MNʲ��r'j	Ҏ����Y+���FNo�9��ֺ����lQ�eN��N�.d�ȔTC�abI�q�b���DԆ7�c\6֚����^�̬Bg�b]�������,̄�^���O�QjY��KKŌڇHU�K�� �4����im��èǏ�h�Q����kɎT28S�=��Jy��ј�F%A�Ha+��
I#i�y��DZP4�3����RU,yF���� t�
9a���������>��w�ӳ��]a�>L�T�&*��P��۟���Q����]�=h�@Ӣ�n�~�@-_��,�"`5�B��؏d�2ڲl[�|�Q�j
�#-�� _�����؁^ ��]�l���!�����p�T��j����Dq]��:4�YŕXl�u���#E��5�w�ݓχ)Z#���2򇠀������	Z��J�9�?�[=��V�w�@3*���aP�? 2�	�A�j0j�L�Ig�U"(d���[$<"9E}:�;�R&�)D� �]�}��w�-sU`2�3Ʃ �'�3���bsw`��uO����1q��G8ϒʓY���[R���G��J�?ouS���b�ۚ+.��P���5�h��DY����F_);��r��G,�!m��DϧjP\+�v4����P��R�[OMR�c���e?@>��:��6b}S�gC��lR���#��q�s��$��=;�^��P���Q]ğ%����v���U38��b�E� "�7�j�+�q.h��^h�x�1�3�z����_F\zT�=>��� ��u��L7�:�����F�C�r�}�Q�ذ�I�	e^|��y����C�_q/�k�j��o������jvf�f�?�YR��uZ��B!��`M���ۀ�a��n��r��W��8@�Lr�ԯ9ݟ�Ȓ�)��:��I�:7��䨵�W��H�rj�8L�xH9��($X�Lm��X�����|��r���Huɋ����C�p۔�^�tdc]��)�^tH 7���u�h����8��$�838y#�o�s�]|�j�_�Ƃ�T+���r������Js���=0�_�e�X�r���s�ȂQ���*�@*����_��B@����Ű_!辩�w��L����|wYJ��?�Z��5K'��j�Z�5`�c�D�)q|�$G(������rR��'ݻX�� �����o�,_�z�m7��\hwpp�0��4;�M�>�i������;��1!s��v�7�ҡ�u���Jg�2y0��|��n{����,D���J�:��}W�$����qg�`G�'����!��Ur��zH� W��M�����=ť(Ƨ���ݴä����51������A{�͜[՝�CFw�6�i�>]�ꤢp8eJ��'Q@A?/}� F���F�7("�9r]V����� ���P���0(��7��7�{�T��DXԆ��۠4Rz&� D稶v�7���S�J��y�=m��y�^��ҺU�Z̭�
ZЕ�җ���~�=Hz?�^���=�1�m�D�2��G"EL�W��C��m�m*�N���D�a�!K����!���*ur^+=�S��6��:nӒt+��Hx����§����HZ�s���J�4�Rbz�tn^-�=� ��kݴ�l�J�3�5���j��I���C�V�j�4<E�n��#�c�u�=�`�����}�'ԗ�j0i�Y�b�qL*� I��/R�M��>iК�W-�WR1 �ذ��Q��]h��t����{��{)�#m�� o=0��ASI���8G��j��ۆiO�8���EVԂX�(����|%��|�{�
�d� �u)�Y��I�$�z�Noq~�ݰ��AGw�h}Hn[�ɋ},c����L��7Z��Cr�Y�[@����u���;��V�����	r6����B�W�1���z��lz��9� U�|����U��p�Pv.n�c��t�)\�/&����RVRz��%���8L��UePGP�uBg���Y	Vl�	����ڶ�X�|��C�mB���������x5X� I�-o�z�%w�T�0��`�k���B��	OaM!��*e:��:��I㌠��e4�f�,M]�IL�/l\?*��ߌ��f��⓹������~M�:����� ���o��Hoz�e��\�a�;��*&Ǳ�R�hT|ݜ�����F2�E4}��o��I����&x~���cް1��JF����X{�u.��(������ay�MT�7��A��ޔ�υ�����UP������2�Hͷ�כ�4���~X�u�l���+�-�g>��R tΣUZF����}���+�v���F�4%d� ���9��z�ґ<��w�����W ϥ�2/{�Q����/�^C�N��U�7[���d� �C��H���`ï��� I������?�OPN�/	
LB� �
c`��#�Z�PF��s=���!��n����2^?�A�!���#*ȨD���o��ś!�E�.���{ 5�hV����_A�;���.�]{��e
�X��긇�^�\�302���>{Jd2�A٢2N�/�oz�>�.ĬQ�%Ǧ����R�Yؿ�LM,�F|k�n��BW��N�"�Z<$� gg��	ͧ��?8<������ eD��$�^�p�P�*�Wڸ���.��bF#�#��0йo؃_�����>$��� ��%Z�^��}�oLy���$��H)�i�U��������@ljt�
Q�ߌ�)zq���N&b��=`����bxY�{��Q�Rz�#'/�B�-<|u;5�=�w2�J����T%�>�<�k�3|�筐[��d�೫��Ht�ԅ|����Z�D��o7�͆v� C�����jS|���7/�����=pB0m�wbuЮv�L�T�!��ҌbVB�BX��w��Kܲ?�o���*�ZӢ��O�4����:��cw]9� r�u~�#,�-��vr�$m�V%�pT�C�)M�@��u����tAF�o�i�jV��Y��%ѹi�b�cV��%j_��
�"^��x5_h�M)���K�3��� ��3�4��1����^ܩ��b�+��\��Ц����n��D���8�#�ޔ�D�-'��[Fy�<z�e9
���f�f�2/�X ��~j?��!�{�l���&��DM�����ύ������n�Ó�ޣW��'	U�yIP��~��j?a&�y��<9�I�����01�rh�&2˄�O��m|/���?����uGB��yШN�gxy�t��!��j���?:������|/t$��Y+)?��(��3� i7��b�#�����ж
�&Z!�th�@�	��b��(=� H�f�#?K9/*E^Þ�������?('{U��w�T��j!A'i� ,�g^�Ak�P(/���r����0є��y�LAȣ͢�c ����Ӯ��~7f�<^�O�?����Dށb�EX�I��3�-�?�c��]Z�a��E�m(�ج�O�εy��<Ч��C����G��W��j.)�L��W8��D*���zQ���ŏJ߱��������(�6
�'��G6"��[7턖wen��&�\aLE�Q��<+Vƽ �����>nCk�$�O�cQ �����1�`��*�ʖ����34fk.@�ý�D�Z�Ǝ]Ь��N�Nn2+�r���)��wŲ�}F��o���	{И��D	�)��0~R�Ƚ �]�v;%��w���
D�F�=�
a��,z�K�����aQ��3*��e�2�o�V�F<smq�N)Y�U�±N�\�22;�0�c��Ӳ��Un����wNC�f:!��
��9'����g.Mi�Z�-.����E^�3��˷cA{/�V,v]׷M���d���mZ`��w���6@?&H�D�i��F��^d��1�9r�`'�ᡏ�<]$�'��no��+=}ˢ!M�����y��â��yD�T�>���l#�9A���į.!#{��n	�{W���<��6O�D�s;hTc����6���B���9�q~$w^����Xu0]�8��#��b�;��:��d����"4�>ݻ�43V���A;#�O��~yC�%���C0X3���Ε�p��HGa����p0JXA���ԊO��yHʡ�2��բ�~�əS��z,���J�15���HNd������ɓ۱M��%�uT`����;:Gu�"�����i;�VN�`Lj1rn�h��y�tw�Z�-���N+V֊��R�^����r��G)55^����>���+1�<n��W���u���mIְ�.�zZ�q���n]�N-����f�=s���yzY^���~V0K)�J7ɹ^�����R�WL���A֫xf��a��*7(~mɈ��^f�K:2�RP^�4u����8���������/$��hR��ۢ`�[H����"rc/24��o���U �)������1t*�T@%��W���U�N� I��+?�%�+L�vDQ>�I9?[/�ф�o�Α͉,L���L�&c�~L���맥*�������f�s��j��(B*wH�ZS���v�_p`N���SkK���%n��Wkwcđ^W#��<���R�^�z2ds�}�}�ް�����!��-��뾍���	8.�V��7�cӾ�ͨ6G��n�H9C��E��]���e��q�@������@(���NF�i��2@{�dV�-��:��B�K�$C��$$�H-ЗA��V�䛨u��w�zS��?�ɬh��ᙂ������ȩa��'���8-ݨ����E�g��8�����!B����摻�AD������Zr@�ݭN'H��[r�*�!��-ަ�:�W�-����M>L��,�>��b�~A䘁��0��u{���j�Z V�����5�m��[�'R49�l��!싚ߐ����t3p���7扇�W�Υ<Ak��L�Ψ4�����@�/\��m��y�	���ȭ3q$�R�n���m�K<�M�V�`���q9ܖ��Y�c�c��˹Q�Dً0[��#��}CAMh2{p�B$�$�f�b�smU��1K��/�ްF����LÉ� J8����Q��8Dc葰<)�"��%���oe�
;�5�&�zv��װ�P�i6���O�kC����C�8R�k-��C��B*?X�N\G��Tn*��?'pX3Zy��(����+]�.Lы�ն�t��ɡ���t/t��þ��FN>���[���;z5Mϑ�w���,w�x��� Z�
a�6IRm6"�����y,��+)D�N�F�����A'K" 6��7%�=U�Ƹ^�`�p��W�>Ef�ԝz|w��.�U@k��1�TLns4I�2�_���ul�e;�VY�\$��(���_��5頋\&���d�+k>_�7�k�~�冠��/�ɰ45.K��m��[Ҵb�X�4VR��w�x����L�rV7c�y͵W �	9�Pt#^A�l�jd��̚8�F�t��z��*w��]��o�Rj�B`5����^+~+�73d�<ot��\NC����F��LX���,.Q��)� p-;	A�H|�}FhG4��}7�/�� 8��FNpʳ�6iLE �l':ݭ����C+�����V"�I��XN2��j8~�V?*����)��#�2�G�sG�����+ox���@���R�4�&%��V��6���m?� ��oe s��@:������6g��"���&Co��9�QԶ���H{'�z��%cG�<�v��0G�Zb�����C|���7q�4� �:�K�T�j��7�?�~��7�$I�F�.���9���x�ؿ��?}�ö�#kgQ~j��G�q��e��9�[7��
���j�J3��-R�:�K~0k8|�������T?��9����t��2����	��B#���u<�zQ#�����Jڼ��QR��bi�o��������1b���X��.�*�59�B3!y7]�0�/	h��#e�}���n��
_k�7�{U�O�c#��ȊU��'Fp7K�SP"0\�\肺츐�y	�(�~ЩI,�A]Q.7M�o6зON'���eu���!No�垷E��{��&Tѹ=�2���v�L�e(���EH�0���+hE���bCy<n�l����}~����6I
�A��^#�t��f��T�a���$9���@��LM�z��M�}�H�N���-CSMM��Vm�+x3���L�h��9%b�k|�`
R�#��h_��g��^Ʃ�A��_���M�8�ʅ��Ț/�V��7C.�4��{�V'��Ԃ�n#Қ�M��DT�En�uB/g�e�F��������l��vςk�|m�a��Z\u��O�s��.Im�A�N�"Wp�c��{��<�2i��R�5�X��.��r	�Һ��~M�ߝ9�=��o�1ĵ��Co��B�1R��H�1�Z>�G�:*�3�u��)���K腁<TIV|�����i���q�� �W�3,ͧ%"WD��:2�5=���?7~.6��DAp��	��;�F&n����Z~W=z�2#�>j ���-�Se���ܭ ��i���%�����9�C�a53���E�~�d��Ժn4v���9�fѮum{"%���S0@d9!���-%�2ߛ���\�Pp{�:��jt�Q�^��XMA$�Y(J���as��1|;&�� `�������_����0~v-��-[��_�����a���z�g�!��,� >�Q�D��=V����-����̜@�[(�ޏdx񈳁������0�}�	�S��b����[�QG6�$JKJ��᫬��+)�`Hǂ�v�u�f�[�7"�
)>1���)p���a��v�=g���6j��gYIe���b�
؞�3�ګ��n�x�"C�*X���<��.��]��ؚ�C�� d �j��d݂��5۽�' �V�UK6D���9Q���&��I�Y���S+=T�D�\`��Q��߰��h���"{�6y<��:)���,(���H��ryL��V���7�d���f��'�H�~(隟<�A[����O��K� ����ՠf�k��a���o��%W��75:�#�N�����0ۜ����7���o��v�*H��U����e�Ak�e/�v?�95�y��f�7Lj)��)�N����J����\��%L��c 6�p�J%DA}o��_-���%e=\{|]^m+�*1!��2����a�1m�����G�O�FO
[�0��Њ���{:͋O�r�P�$���$S��R[�20
�+q8�wD����5��|!:�<��囋�	=�����	��Mö�����4�M�:�(�!`���8!��X�'��9�r�PyJ��!2�p�*R��� �Ѕ�/�s�2�8��߄�M���^ʷ2_�xb?�԰HY�{!��n����}�
Y��JAP�Y�R���Q�u>��!��܅�n�����M��4���
E�|e�`��A��ǛqW�rBԨ$1����j���4��$��ɡ8��7?�hW���n����}��&�v�1Z��z�  /�]8��Ui�˵�!r@�@��G`��Z+IKa����8�2:0���z5�x�J�O��$���nn�0T{��v`�V@9wN_�'_�^#A����V�Uc���kLNh�� �nKabƑ@��8_b�ː��	-�Sbi�S��f��V��$oS�پ���F��o̓Wf���)4*�i��o3F��kbF�߷��������w��B�������ֳ������yؔ]��U����#�֧
i��I}G�+6E�z�C�b��3T�ٔ�����f.�I�m<���$rǊs�Iɝ�2s��Bˎ=�V�v������> %0@e���UL�Z���w(�i��C��{]���1�&�o{�.(^��wx�qJ�n����E�#6�@y�h%�b��z�*��zw8��=��O��q�ͣ�L�oA�u�����(�~k~�kV� )��3^�����s čtJ�;���+"$�'�PĬ�}��ğ��Y���g�?`�I�������;��io�K���!��xh�07-���ە�*N+}�oW6�R�w�$�wg�� `�?�|�؞r8�tf���*GѠ4xaf��Z�u����cGZ��Yu=�:z�$2Ҋ�`N,�����r��=Z��z�d�j���<G?I��[���p%I��Z~�ī�(��_�Ȣ �d+�#Z�e�_���i�1��GJ�;��mr`E,�>_�3���n���Z^��<pV�qϞ���{b��4�e �`�+�x�O�0=y�l�oM�u��JgL��@Fr�O�Z\(�怗�o2��=�9n��o� {w��8�� G~�o]I2�S�-�s��f}XW�>ǝ�

�K�Z�=H��@�7m4c���C<���J�1+7�n{���r6�
Vjmx��֙�����W'E����C�f��䊶2�f�&�4�aS:�$��p�Ph��lv����!h���֍�=!Ab��Q;<�����o�s�l�Ǐ��ˤ7"�� \�,PF�)�=l��f�!X,��J�����煆�7��LVK��fh,���#Hs�0+��JVG�Oݗc���'��Y�"K;R@�A2ږҦ�$!Xg
��4�;��ARz=,���EBuAk�;Zk��C?N�l�H�)\hᤝ�����F���$?cL���=r_]��>>pk]���z�b}�D-���*b�=xo�qmF&�p�z�עc����Bs��<�Y{�{p���~Zuh�(�F�-���e!e��O����p��ux�<��W�`�.�3����^�����u,�QE�r��P�?����+$R_�OuH��Yo��̨4Ac�g��m쫯��4iL���iw�;i;�$h���6He;��w��(�V�W=�\`n&55�y��Nŵ�c����'ޗð�p�'�_��'�=E�����.�)&�`���&f~���=�����TF�{�5���<l�\��lX�b�o��^�
�M��x�dW�� r���{Y�OC�=�cb�������XG����:a"�����w�x���������|�\N�曅� �?�2�j�7i�Q����"ؽ�3J���?�������y�ؼ��R�2;������B4�׉�j�1���Ɵ|�$�������'��2�Y�|�Ú7x ��̑*�L��gZAv�)�7��� T��Ux\�q2�՞�B,N-� +.)����x�p|,�����~:3G�Pɳ�?"_�$Q�@�e�e�)�}�I��,=����F��Y��/&Gp��o`!���4w���{%$s�ߜ1PY��z��D�,ֈ���*�w&/�픥�B��q\v�D��~�l�O.۽�91U�	�lJ��CƫT`��Я��4���l�,� C��/���e1��W3G*%}yn5,��-�m!���Lmt���lM[kY��%ą�鎤1w��@(Q�S�u�L����#(l�W��d���X���FԮ�f[�a�fρ�:��Grz��������$Ī�E���6;�k�oq��2����آ��GOXT�s��%����"�TȈEC�۬T�.%�R�y��B�c��%FJ�k���W:'݅/6<�G
Ƨ0�Z������bI<�7茿o��g;�	?��:or4mπk�������, ����ꛣ�(�����FO�BQ���3�a|����hg�ݺ�&r8w*�%����hL�,N����씅���`�z�E�(>Ǿ�N�eG��^��G%/$��[��U䡢�}z�tQ^�b#X:�n��u���&��0j�T1\�DPf�`�Rm��w]���8���,�Su?H���.��K}hu� ���:H���h��?��9/e��U���op8!��f�?�����Ԟ`���傅Z����X����&'�l˼B�A̵��&���'I��̮B�m]!/W�� ���N�����-�=�MW�E�s�$'}���"q!=�L�$s�jW� P2��^�Q9�M{�U)����`9��D)7���Q&��ݻ�EY��>R73��le�����ȥ��"�J�,�Ż���FVJ����'�~E�y�X����Y�ث0Ź��E��
mP��\�%x����8EG�CKi�87 \��~�v{�;1�+��b$��]���ǂV4Zo��@��~߅���B�b�r��X� -jB��������(��C�֟I�o_����k��ȢN�Y�d}�W�����M*o�@XS� ��hYx|�����&���6:�c���jT�4��xR\%�~�
�#��k��LT����0#�İU��I�׾�e��EzP�����5��d�_�E�1���{	�vw��ѻ��tFm+�K�+^O`���� ��U���g�ͫZQ�Xþ3�Gi���p�:-���&�	[�L�,���t�(E���G?i��Vt�C/0�-"���L��|Fuo�l���n8�U�ʳ�C�j�C�l����;��`�y�d��2��}.��Y�,s�iZ��s�.���Vr9�W"��a㢌��Gjm��G��٭}��~4��:�LU.Z�2 b�U�ߝ"�f�<������j&���M_���oO譽kVA�ӶFO�1�"D2oH\��%г�N\3���Y@��Lc��N�?�6ݭe`�3ۦU��kq�q��+�k��_.7��M�>[���⛄T_�軰M�D�e�̡	ck���_�4U�ڜ�:P���V:S"�;�3fA�<������@�U�#��,��5��,~�n��H�p����8�κ��e���C�H�s��#�B#�鈐��?��׌a}iM��M�l��υ�6��+N�ǣН+�JLP�(8z"�?SuWd��tms��i�^Vh�C�3f/�� 7x	���f�*J{%)��yJ_�I$�a�+�x��EC��F�"��̢��v+bb�<!s�ǝ�$VUҽ��j��bhp��D��4}�m���i@�涡G<�H�P���:��%�CǛ�gS�2�M����IH��M"�y�<�I#�V!��J	�O�E�yNu�l�1���K$ԁ���({���<B������%��1�)�T��01Ɵ�U0T$)�B9f}����;Ui�t	��ℼ; X矱���
���Вj�e)ZO�]��-�.R~a����s����O����*?R�c^ʡ�; ����w��↚p�-�>�k��, *������
��NHPn�W��U�J�9V�e9��p�s�ړ�H����יx��)O�@��\�.ݢg��K�ȏ�J�Uk�hg�#y+���w�?�F�;@�Rܐc\��砺ã���t�G=["Pޗ���5u�sq�T�5��(`�r���![Ri��_���RsM �/]�r���6@ϸF��y픔�T����9�SO��z�E�H'}r��f���Vh�!$1SnrG>�
�X�\���t��cAI#�.QVӡ������
�?�BS0�yEwdg�e�]�lY!`��\]n�EseUy��j9-��p~x�F��}��і�* :
�����p��� `�=��,r��-D%;"G��0����諸�"��K��bĂ៳��#sɍ��þ�=��vD�)����칏��r�W�eUp����fNN�;S��~i�s��4񫓧���QE��fiZ_3GC�X�|�ڪТ�"��7�ujY�w���7xdo��%77�v���� �\0%�����Y�a���q��18wڠO\��fu�n�_u�{���2�� �~�N�/���E�]��V���{��K�DEJ���e��5>v~G�D��>{[�g e��&��/za�V���
�}D�ˡ�@R��v4�(%����b�;^ Bt�tȜ�7B^{4�q=�Yx�v��A�˧��-�bφ���"����ߜ�o��E��{݊!�J��A�kW��_>�4H:�&VAm�/��������S�2�p?��ׯ}��1�
T���sQ�b/YS*���R�V߻�+lh�bAĖ�Y/H}��r�w֐.�]���=^�ٷ��$�9&�]�I��B���!߼�j��jʿ��l$i�^��<�z�W�]��j[e���ݲ!Lw!�'\�ʭ3� �~�#ܴ���-��`���:Z�A@�In@@�'�(������ZG;���K?d�'ٙݧ�ڃ1_,g֓����&Fvw4�aBs�|f\�p�;��3���u�^v�s+-.�V�o�u��@Z�]|+�As�UU����	���{�����J�^]��_08�l��:!�n���yZ�v�3'�����8�s��-�։�<FNch,�y !S��ne������`����uY�@��M�o�2��1������E΅�ե��L�����A���R��ǧ|�c试���Ҿ�r{�!
k'�U-N�
#�x(�Ds)���w�����2�&�W��
eVȸ^&ECo��
�YIq?��՛7M��K�`H(���'���AX(�1s�P��=̂�y�?�gE��v��U����+7�Af��Z#��:�C9<۪�C ��Շ�X~��KZ�pv�k�ą�������ny��(-��>fG���8�bj�~���!���7�2K��t�SȵM҅����C,��!E��궬����F��	j3�"vas���T��d�¥y�]��K���W�"<��v1LB,��h��O�-N�N��;���s�M|"T|�5���{�AI����bw8�b�rv>�m���^�4��]���	�#o\�6��xP�zCˇQ]������Yv_EI��J#�S�ED�a��"N.����p_�`~�z�Γ�N2>����wr)�I���ޙ����,',��HǙr�����=>+�"bM.��-|�P���A�0�+�c�mEC����2IM5�Q����,;�?�{���B
,+�b�y]�i��	9Y߰�0ɖAD��Gk:�����	���� f�,�
�{��^O$�P�x����?�����6�	B�`�@��:�Ja�{�I[��u�:�N<k.�b\H`�>��no���[�T���8���:��CO� �\��<���2�Aǩkf�M'^�r
�qU2>�MG�Ġ/�������qP��z>�����<�u��F\����U$����Q�0ཱུ�)I�/v<�N��l�P�����u3�k<I����	HB��n*��^���U�:2�E�	�J�34�&<��fb�m�j�t8q`���g��Ar��j:ۀ~�8\��j��3�y��@�>�;�G*W��JRya��I8^�t7��Ҿ+HO#ֳ�1������7�l���5xL��gC`sM�H�&�<�2L!����������|��4��w;��Ϩ�)]�j�d�#�ب9�1����q�<ddؓ��9� �ƚ����9
���g������З}��Bld��Y|���>��餛��݇�b��iT���~=X���W��K�ŷ��J�Fɩ3��qe���ӡڎ�ć���'V6�20s����J%��ݶ1�^{u��9�[0C����e��B,���a�Z��� A�n瑦�{�he�L���@K�O<�G������|K� 3�z:���9�wQev�C	�:�L��_� h�����h��\~�\�rY�<
��GU���>2D*�T�GO�/�K��,yH����;q�I��:����<�=y�/�{�^��
�Z!r���������,�� M�5CpJO�~��k��;�շ�\��X���jX����].�a�F�l� ����L㿾դO+@��@Ȕ��sH}nw�t�o_�Y�^`%_����lɄb�/e�Y��=�l�$9��[�~��Zħ��{�ou�^2�ߋ����~�k���ɝ�I��F*��b��k'�e����20X��f�#��^t�y?��;�ł�	;r]
�n�e����W�xJ�ee�&�����֚���CE̺V���c�f�l�[��7�)x�^��,N�P�Ĵ�'Z����T�7�c9ge��-\:-��U�:�%ۭ����\��>�`���pڥ=0Lj��7����M�Հ�4ŀD��6}���-�M��N�gw��f��Č�UL�4�+�O�v���;&�1����_���\�ЂH�M�n�[c�]R\��V�<]K4G��&z��:��\h|���������ߪ~�Ȭ�po!�s�B:,���L������LS�Q�Mcl�r���ƈ8a��1�@�����G�*a�c���@N�V�� �]�������va��d�R��E�+����i¹�R�	R ��GU2_�� )h�n�w�h칥
kZ�y	~�^�dn�\4�u�| ��÷���� �}O�s������Q�זQ͵�[n�FqD,�'aj�r��)d�����!��lA�	c���&Uֵ����+�t�X�j�0��Kw��u�rJ==�aVM)H�m��p,B��@�
W���>��(���Z\h##���z���v=�?-��Ϯa��W �
�@4� 8x/yRl��y_m���\I�p 8���(�	F����;���s�����X9k�N�BiՕ�|p��04I�s�:	a�*��-�}o��Ь�X���%��0������M�=J�U�*Ʃe8�hnё�mȼ��՗������-O���?����%�^2bt.��tϰ𥤶�Y8X$n[��G���"&��ʞ ǈ�pnYh�C
^ٍp6��Ӈ�/�����v][KmG�[hU�9j�����\gm��~Cn�2q8���-4{�T�@��aW���kzk�A�`8��&�*�o�k��ӣ��A υW׻�&�2B��(E�`��������XAH��F��8B[�Ӊ�v2w�R[<Ua���d-;��q#�g*`&�Y��3�/�</���#Qrˡ؜��������/ԸnL�v��	Q��������>i93� kE�"��?�k�,D�Q!堭�<��f'��W�۴�^�5��v�����,+��E������Ot�c�����j��E]BK��g��	9�0��Id�����(�<H/��+)8���#��(��'�y9V�^�
3^[z|zSb�+�?�,}ԥJ+P���s���trl*��پ,�]Y:[_ ;�~����h�U�t���!���3ЍGT�nם��N��F�K��
n	�mɩ�f�vȎ��+5�<Z�Uq*��������/�h���)u�*�\Y,B�tPV7�v���6J��O���j���x�һ0a�K�Az����3��0���g�*���P�I��j�Hѱ*<L�.�;|_��M�oa�_n�����|��._���0�*�`�˜��D����څ6	c���T�nI�dgm��V����1�ݤb-���s��)�j藄z%'$=3����J}��*�Fj�o��3�z^��gWAh�\(g��ZN��G�9˨�'I �ja��4ꄲ�C�^����~ܢ�}�ۅ.�JjeQ��6�c7���Q�����wˉ�{��8���MdH�����8B�y�Gn�rJ�7�D�9e�6z��Z_��S����&ʹ��׼�xvE/R� �O��Ϸ	Ϸ����hg�CSy,���Z '$D���F��z9njr�����Lt��^�k�� �Z�SЪ�6nv���:�2Gm��h۟8�0���LYh�ϖ������H G���yGoHV�,�v�\B2�x�����ֻɖ�֡�,��0��Tcy�Ė����wُ�&^������d&���YL&��m���`ʔ�I��Ea
Oz�?p/!䛩�i��V�5���y�P,�tw��ו����%�H��f�M̽�m�d��XI�nBi	�c=]R��d��"�fω�̕y��*e���1})�B�8�3����eMA�<+�>�47�_�e���Q�i
���us;� /��V�����p,�r3_	�C0*w�A^5�g��#]9��9{��������5�ԼV�p�m���j��f/L��@�9m�+̚X��o��Ic����/+t����k���|"R���������`�����r�G>�m�QD��VH���Y�귒�ձ�P��j�~U����/�fN+��J4@�6=��@����.�^_���F7-��tAB���̹�i�B�7
!�@o&�ڭp�T���i�˵�j��5���������'�{��P��,m���_K`��x@�;<��]p�fV�
���;�'���хDO��mľ�t��$�6J���/L4s���L�������[B�z�=�@�6�I
���f{D�=�:2�F��>0�<���X��f����J:�1ăJ�e��iM���:ᰈÄ�:Cْ�S��+�R��~,d�I(����aV u+�ae��z����.�=�ҧ��W�����Q&7-uU���
pOZ��Ȧ`îq�~�R����IEx��|$���F/`w%����em!�q��7�bFa���።ܣ,ҟO�X� �^���1Q��p]!�|(���a0p�PE2NMX5{%�3�7[F
q�R�羌�DE����2:u�]�G�����!k첎t>�C;
;	ZH��b�Jt�UƉ�v.�>�<��A�C��Y�X<}����<D��OIOǱ�> �d'�ʃ�4K>�3A��$�TN�2s`�1Hba���L9�$�yB/��y��ԋW�0���f�u�y�"�#b�t�q{k�s1>�g������Aj+�na���`��\I}s|7����3|��>�R�U�w#
ᵕ�FԶm��S�د2f�Z���3��k�?��͞OWѿR[�{�J ���,
��o��=�pE�c9U%a�u����y�G~t� m�>p���p_1�w׮���gv�䞽-u]n?�3���{p�g�Kc ��|S�[(�D���6��.�����-��v�]G3��'j+��\��z�9N݀�7Ʒm�kiA�����8����?Zy����'O��k�-M�Mn�{��ʉ?Į;ֹ P��U?.%��-_�_!��x'��0�J�YE��n�1�Y%��.�evC`���ICڷ-�p���%�o/��x� SA���j���	�E�l���I��\���J>�1��1rn�`�㵨'�	e��3&�a{6�:�G��Jx)�$�����i"#�_'CHU��@��R"P
�r��;uo��4?�o�0r?���΃��	Y��������%r� ͬL`�L�g�X9<�P/�0t񻢐 2����h��֣`۬��~%�>It�c��6��R��]��$�of��s��Y���D� �>��An���Z��?�cJ>&�c���SK��'`�\��<����8��i��PG,��]��vU�\���M�̠,�q�h���g�l��0NB��`���9Xt�`���0�.O)�-*�ł�_����"�k򛅫YDcr=�t��:s���/�z�SQi�-~��O4�����qŌ���(6��a��iG_S�/��W:�'�B��o�^�5B2*sS�n/l�(W�]g���=�ɉ�Ge�`����;n�V��M� �A�}"��%mBN�L�
aof���~���V]��!�d��f��[�z�X�>i���#���L��*����Ǩ�Q���T���0i�����7��[5=`)�~��bFn<����<�X��հj��pW���C��X�9@_�1����nc戭(2������i&"��D��e�=����B��>�9�i5��	s�_�d��� Y����Ar���rkEpn(qx���Y^�oI�=��� �p@ҶF�%�<C���&���,�#Z��.E����U1���#%�R�of��e�]��n���糰� �
�\E.k�uR_�m&�|}���/#.�Ix"�9��E��[p=��z�"1��ہ�|�N߯��<��rQvQ��_�L숫� y�?�z���Z1�U&�uS�����-��Elp���m���B}��+������a��S��aq�(@`5)b�?��8�1��I�]�F��cw��+��$l����~���+"�D������2�"��J׹S)�9^�*����k+`��3��L�Y�k��깆� ��d���~�,��e�"Ť`H6��Hd� ������pi�i�����r��U)Q��pD�_�rd���c�b���s0RR/ՈI�i*>������^z'�#�VC|��M{uR�����V�<++���D0sz��r�"��j�<��=0�+;=���P�tQ�u<�s0O[w�k�Hv~ݰSm�(L�~�4�̎�S�0�w��|��f}q��V���/����]"�pc<����t���ٌ�/�8J����ʣs�ۉ�(�_� � ��CR�'�m��U\�Ԋpـ�Q�	C,�\�u�w�X�YT��2+x�tcN-��G��#.�$3|M���O��x�M؉]VŬP�|����Bi��Ya����O�:�Q����'�ݶ^���r�H��M?G�P�l���e��ǣo��I��[ޓ�%����tݵG�!�Ö�]�l_d�-t��ً>�]{�0��չ�94�b�
���=`$��i3����
��:)@���mQt�l_���K
r7��QFt'�F3�݇������ҟ�6埣����2';����K���J�|j�`�V�b;Oe:���<lk��w��TZYܺE,�Qp�I��}������R�_elK��@�;�a�"-2|���.�Nm)
�ǃ����b��B�]�^2S�]]�FB�1���Q(���MIxL[�6��G
1v�>	���>D#��.F�\#*|nj���c���e�����ތ
��W�'�tǼt��gޜ�1Y�Y�T�L���2��aBV�H'yBK��W��I�{�H�����m�[����H��|�xB<���\7���ىW����x�/P��� �w+��V�Z��L�8`C1 ˟EkASq�	;�"vYFhS�<��#��W����D�ͩ�	X�u�U�"%I;��'}"cM��5��]��l�[.�w��+��o��w}^h��3`�Vl�V�|0A_��Sz?�k@�h�h�bñn1��$9���G*���s3ޑcQ�œ@�+�-�}�� BT�Hh&���`�o�pN�l�N�%����Ɍ�4S�±^��F:���{X%`�變�܄N�/�<4�8��Y��Fτh�6�H0͊Gi���z�7 �M��}`�o�`0��f�HQ~i�`�;y�f�-�-4b�,�	[��b��&�I���f����q	5~N^�Z��9ź�Ycұ����&Aǁd3�Hj�o���M��W��<<{�dL��6��KtFA���īk���*�l_�p�)Y�\�����?л�v��gj�ý_����剉����9kV����\�p��01�]M}���>^����U�϶�>a���[O�����\:�zwф��M���2O���#d�Yf.ƃ��"jM�+�I&�� msӿ��@7��5���\����+�<��1�Bi�� �Y�c-Q�ai��|T��8�%�M��W;/R{�Z]LV)�Er�S}u�ӵO��l���4E�D�9��j�K	�	�`0�
�/.E�o�{8h~ER@Q��*��%ʜ��\�l>ʺ�5C姸�K��ͽO��#vW�{�"Za�uTT�El5ڊ�����Pݡ0���	��� G�w��f�
�,�����nΌ�*�\Uq[)�to&���;n�"�_!x����V}ݎ#Ĝ
d�{�@^�v7��<�^����8+N k�5,'X�Uu[R���煝�h�6��,nYkk�+���&�؛�T\���ؼ�Y��F+ܶ47�&~S�F����MM�B�V2�:޶�e���͒���ͳ�`\��Q���g3�u:q�ꂓ�f���ο��th,�� [o�8 ty1�"���+�J~�SN�ϡoeM��T�n�aB��!}dp�8��YI��S�X`	�'eYc�q��{dB��T��X�����|kJ�0�j�����4�����H�ͺ�"=j�#u�����$���� �~�>�u�&�	fUd��������� sd�M�*�E���G:�)����qf@��J-Ɖ��k��\[uMM���]��Dif
�����,��K�}�DQF���H�yc�_�g��q�<�p�^�N�B�-��hR],��3E��J�N�B\f↡����a�68ԉ/p5Y;fd��N�f����O}fUe�k���C)R�tH��h����2���N(���cܴӐ�U=���>Q���S�:�/h���Ȉ�����5�У��@P �!٢lt��ٯ0�^b���X���S�_U���1�&R�8��e-J�Y��_.������;�3/l8�-Qˀ8�V� ����u~�d2��\?T<�m�\b�]�ǥ�4�H��ѯ�u�m��r�>q7� 5�0�٦���N�g,�B��G��?��F�oB���?�*�郄Ԣ���Y&�����{Q�{,k�]�QS�g�ۖo��a���@��ɿ*�R-������y�<cL��/b�zÞ�w��t-�¾�F�;~&����Sz+*"���ݛ�<檢u�|�����"m�[�nvB1/�������ȱ%E��I�kdM.������bb���=x_~&����Sa� ��@��q[��-4�4�	]�K�R�Q�Ǌ,�'� �=��ǰ���t�߲�}�Q�ڹm�K�}A����&�5�X�)ʁb7�������j�����58�9$��!��j�����e���!廲���QQ��)G~٥�����!��ic$����R%��F��`�sG��Q�,���"�b�o��`��Ӣ���G�a43��.:��ɴ�Х�Q�Ż��Z1�N�=���A�Ҋ�%�ޑI�|;�QI..YW[o���c*����ғ�7�߁��:��nk����[���x��?c�d�B%��qy	�7W�������5N�|��&�-����e	9�s�g���b�E3�Y!>6��ﲱf2KHS��W|�Yv�Sk�nҔY��Ӄ	�7AT�)��n*�p$�t�dMn�X��QЫ2����[	�Yɪ�V�c�2��0k�XU&�,m����lP'�KF�F��â�69�ˣ��9O��#����g՚���2el�| ������$T��v�RE�p6���@@AC�s��7�X��� _�ʱ�C$��w
֎�f�/��}��Ik��^��șLx{��ӗ�虳���F�`������F�0�
O��)�D�&��TpZ��2to��b5M�n�>&�������>]�LQ�׆�g�e�g_6ۊ��4L]��J@_�3߯M��l$["�����Qq���-c�t)��8�"�>P���u� �̌��՘�+�l�S�T���@8�m�4�����nj���#�P�3�h��3��Lde�(�.Å�+G��(߫��������-!���\��W?o��n\��Z�o�%ŋtyJnƄ���5���s{�8�F���r@�m<H�6p�'���hv�Y�x(%�I��W[�뻻�Q�MU��|e���q�ֹ� X���!���w��41���_h�f�ؽ	�w=7�?�9R�jd+#!0Q��Ab�H��|�#��eeS��J�i%4��*>O&������Py
"*�0>�zA�#쳣�����	�T|ΖU:�7��J����9(f���������H��R˄����fN�(:@�l8 �((�M�Z�-,5(��?�����t>��6C�)�!C_g��e-�1}��H'z�6��������� /�I�D
JUO܍���Z���uF0APy����p�{�!�Y�St����\B�����/��M���NF�ֱ�|,.��V9�$S�%ǋ�D�Q�ʨ��>S<�*|:L����� ��,����
+��ʺ�R/���}�xL��gG����>!&�?ib���LA�L��-�N��ρe��(Z����ሿ4���֍�d�$�8қ{ƤfNW���F��pY����noO�����\��8�����é�Po/w���l�o���)�S���6�ܬ����[���S����0��:T�b��h ��2y�K�y���`|#�I��89m⎆�����ֳy8�C�D�IFR�6&%�$a �B�&���`�W\҃�,��l���I~*ś��6t)��S��
�E�+ku�ڰ�^-���P:u��-6�r
����+$rlE�U��Rܹ=,>��ۼ��)
B]ΒoZ������yR3�-o�����VS&�g�Qǵ��ᛣ��Ҭ��Z�8��'}<O�k��o�a�>���'6ͽ���|q�<�K�[6[�z,�?tl�ӄ�,슚[J�M$EU�]��Mc�׺�T�p��g���j��jf3��h�P�A��Ԥ���0栩�)�g��PF-���t��PU���$�߽oq�]L��+1�L�M�Hx�A��>Xg��(��V�?y��%��0b� ���K�%�!1GJQE
Xa���B����۞�E�a0�(�MY����J���H.�Y��9�s��~	�1>geTx�B\T�����q�t$��|U&��R+�����^����qH�o(�[�	)�� �Z:>z��m�m�z�<]H�������U��qZY��N� B�����Oӧ����Ix\�1̑��'a"ˉ=�j3|@��:���� ghK���\���"�� g.(�A���u�	h	OH��ٖ��G�t��3"�v0��ݹ���|���M[7��ڬ�����Sk	�y~,6�Gg,�(v^��;_�w�v鴁��~Ԗ�џ?[Y�0���NsE>���O�_*�QH(�Q�4'Q��a?l0�#K�a��2��`-�!���J���1u���b6z.���z/�*�\��t L*ja�"����hC�>d���0{��|�E+���$����p�`��.[�U���k�s�f/����ճ��#�c[d���(����T�WE�o�u�a��S�I�YgW���N�S�ۭ�k�]F�Be	��\���L����d��@�H�$*&���@�o^��x}S���w̯Vҗ��� d��_h&�������^_7��U��L��
�ze�$	<��ۃBE������ˢ��ݙ���w��q�n�-W���Հ���ڛ����\d�aO����_�vǷ��M�
�5�[ z��(��?��b�g�Y��%�(�!�K�e�EN�B��]j]�+���REU�8ҵ���&�E�J��9��q�Xx�[g���%��WǠ���鬏��K��3�;}ȇ�l5�P�x}��I�U���` l�ށ��4�nך;�u4��K�gi6Q�̜y8R�1�q~�0p8��ƀd��h��ݣ���6��5��MG��[�"3�ڝ��~�100��Q�I��7��v䑍%˳������GŲ��Y��"Ǵ��;�1��v�INF�9�W�LB�5�k����g���7�G	w���n'{%?���Q[��6x�X�<]~��n|��G�^o���>��?i4����;oE���dY���So��� �r��~�}��= ��k�g�ju��f���ǂ�̪�h"ӽ�M��/pǆ��C��-�2�<h=�d>���Aڂ	C|��������/�� �'��C��}2\� �D�����yF�&E~ү�nq=d��9i�gr"*�\eՃ[&R�1a�g�2��:ʛ�� �S�*�Y
����P�`
���ۑJEL�2�3 t9���g�d��W;O�50bMuIUv�(�ot?���N:�q���z�y��:��C�\q��1޸�[���C4��<�b�ؑ�6�w�Q�E��E����/y��A�Ī�!�vةzP)�K0�@���R���͸N�R(��\63i�7;�f9#����m]w��N�XS�Vy4�(�!.ֆ�!d����v��A;C��'P34��Mлq<���r�&����L��d�R��ul��}`M��2��-��cm?OžD�z�<-��X���Џ�1F�<��Sͬ�����v|��ddH#
_��D@諒S��&/��6i[���Hs�'U�\[1O���[,T>Q�K�#a�@1S˘�*���)��;�H�sr����XyT9��~]�G=R;��.Ӌ�%V�o!I�s
� 6�	�a���1�J�37�"�±��7OΕC�w}󬏯�Bڢ��"�����d��D�Q���Z���l����^ӷ�q{��TU���uk��H�`FM�FC����tƼ逭�<
Ri���[����f��7�(j�秥��/�mt56���N�.�b�O� b[�������Ac��8A��ȝ��R����[�Y�Ĳ��o�x<僑I�/׵Ĭ�0�4�a�dQj��g>��e��y:��Tz���x�$EDY��r��h�Ik��eX���Ӗ�-�^	�퍽�(FUd+�&J�>�"���V�\��<B-��P�U85����Ln6�m[X+�t�ԃ4p��Epѧ�P�#�tz��GL
��-�qWfJ#�N�J�il�0�4����2� [jɞ��7`/(տK�Lik�	۪��,)�]z7�ȉ��Öa_��|932w��Bw��C	(��d�L�U��a������W����;�(ȋ9cY���L&b�P�4��&�Y��z��+��ш�O>���S>��C)�l��Q�)��ȹ��%�{�(��9�Ʋm��X�{����	�n���!� ��j���p����R�%�wڊ�kb g����z�=���Qc�X�_<�K���5�a$�A�b�dԂ����}�#��z�t&h4�J��萛��3L^��\�4xI����Ss.G�*�R���4��uDdQZA�5���Y���؞�Vr�0�s��ë[QxU:E5�_퀏��1 ��t��Nǻ����9���j���6��>�R�K����1NJ��nЈy�)�R��)GE�'�zN��X�u존1	\5<��E���)��}^��e���1p�}�	��a�,��r��IOO���ė�2"pE��m(�	w$p�P��\F}H6�S��<�$9#;];���&S(1��M��LW:���Jk�-Vub���Y��.)�l3jܣr{� 1�ڽl�|"����?��r����,��*�\�԰�)j+to���B�����ٯ��z����P����yDJ9�:��F2!��eW�����ҡ]�c�t�+�٦Յo$�w~�g�g���c��`�@���K��mq���)�*>c���6Q��g(zl��RAC1��S�����A]%9`�4�,���?����F2Z�o�"���^Pӯ���Ÿ�FS�rF�%ŝe���K(��d1�ヂ8e��w
� <�9B��~%�*��DKQ�M��Nk[�e�n+�E^�<Q�����]C񵯁�h�W��5(Aa� �n�I�A�� ��[HΚC�#�C��2�������u=��Agy�Y}����+8�� ��`ƍ�7ⶥI��q��~�U��	�nuڰ�$Gy�|��y�^�w�*�4x��T�������+����i�i�Q�@�ڢ�^Q,�G�5� ��+�1A���� ���	{{f�?�A;Fj����5"�$��U�P
S�O��x���1��T��Ҏ�>�<T����Ip�skCaO�(�&f���,�o�"���£�FK��"��sD�d��k5��CO�*n-cb|���X�b�e�{K����0��f�#��M<F�*���\(�x�pP;'V{�}�z�54��5�����,���o_�L��wT��5���k;�*fm��{OYe�j\�6K��9t���'*�BK�p�ݨ���(���	6S}9�N�1���p���#2���/D��I��b��>����IWµIQ��J�:uݝ'��K��?jj"%�<��x�]���y��50�fὑ���%�7��ּW�쐚uw�9�����7��>ps����z���NM��A^����I&[�x(�s�T�"}u��ѧ�'Cx�`���r��
!	����Ơ�٨'XIb�+/���v�(;c�I;=�yy3P�W��b��0��LX��Qu/�A3��Y� �/D�M�U��ߜ����Qm��:�JU*�`�St�2+t�L��r�%���%e�˚Y��r@�˚~ xe@>�|˿"��>��7�ݪ����F�����r�Cs��=��{98�����Z9��Z�Q@F@)�&��UE̲g����{�@����8Σ㉗Py��Z; `���f(���-�
U7�{�e���>�:+%0 �o����{.eX^W댞v�;������9y�՝�W��@�����L>��w,�.-C��J��u��ÁĂ��J�e{�Y�O f"�Jo��������$���u�7�E햴���� y����@t�M���s[	�\�S�N�4$Lϩ��D~Z��c�C����O��|%��x]b�DvT����y91�EN#�T�Q.ۚp=bYwO������o%��:�&���Bn�L�<)'/��{}�I*�9��5,���7��`�Erj ]�?��yQ둽|�]�8�7���'>h[��5S<9Ի�
&If��)æ�B��d������� ��<�C�4G
�J�Fy�Q�p�֛��$�I��v͉Z�<���Fs҆��E����ؠ9n�8�����~�r�*q�	�_s��2t�ݺ+ܱZg�� ��ѷP1�O>����[=${e3GNE��5�4�"�.�R����K�X7�xn{V�Q��0��,��%��i�G�������RrZ�g���ʟS�f�z���l�A5+��NC"o�g~4�ˆ�ߘ��}��8ڟQ�+���խE�ލ�,0�,�@�;��l�ZP.���ቨ~�����E�(���-���U�/J���঍���A}_+����J��I0������Jq���b��|�dЭ�JV�1���5Ӷ����@Ɛ{�
��I�D�8���%[��={���k��P(��́��,�W#��K�R�)�s1(=��,��Gc����g���AR|�d��tɡ�GCd4
8s�E�����/*W����kʬ}	 �-����H��=��'��7��4!D�Μ��< 2U hho�7�Y��P+|�86��������<���_eh[�g�k�u�w��*�}`��N���|&�n����>!=ޢ�o��j6�/�@��I,�\2��G.V�8���Z�#��JKV�e�����}�?��q�I����n����?,�ħ|�v�g)Y�0�O�����YD�� �ѓ}�5%�Z�����V�͏��tؒ6���8�`j�c`�N���9���5�l6 Q��yU R����I�-k���m�����.Ī�$"-���'V9����
Zݦ��ܗ�?��-���߇�d}�@��1��6,!� �������~�o� h��6V�/�:�q��2s[�ՙC��#�{y�m8R8��_�n�"�>��ś��ݘ�l��49xe.�D�`ƛ ,`)�b��$�1�~�����(T��8XTՒϙ��������m?p#�7i~ ��}��yAPe_�4����0j�r�K�n09c$�F��Ō?)7�O�ǆ=듁)�$FZ����!B�q$���50FH�<>}�ؽ~�&ഺ��	'gW�O���[��rZI�B?`�Z�J�lF4�C��^�M��	�}s�L+�¯.d8��_�������gS·��|d�� ����}:y�վ\S��l9�/IC���K�yU�S�2|�瘺� ���!��J�;�1ʐ�f�yG�ey���sͨ�6�.��Es��{b�\Dݶ�ʭw$K1Y��)YdA��Z�N���� G_2��@�hE����y���تy9JK � &����z�3V>�+�T�-?�=�4�P�&x�2+m.����=�T���w�E�.���ΝLު��i�9�8V��4ͣ�J[�����4q�4)�
G����t�P+t ���(��帰�����&�^'aY��Z�qj��{�ɖ5ShoH�y)4�����P��~<��i-�[
���h��Or�X,�N1���0B����[Lψ�nu\;�Ϭ��X��2�9C�#��:4"t�_F��2m��r��
�J�;��p�(@˃k9��>xt�EMf�g�O+ZAqdgFz��:h�Iב�'�����gE�bY��;Y���?�U_"L��f2����*D�q�o��w'��/����6^b�L���uU"�I>stY�5�Ta�D�P��WX�T��׀0G�'ዓ����z���A�o��`���M�Qk_S��ޙ�C�Y#������jO%�LGUl؋���@�Y����C%-<v�����ε�?�&�6�ڃ3�c�:��|�� ��z�uİ�'S���rXE�Ϗc�o�@�a.�I��A���K
������Bǌ�3�ޒ;Uyswg�����$�����^^o���|'Y��ؤ.�U�>��Q�cqV_�v�U���a^Y���P������]������>x�������J�_�����P:�)�� H���әdl��9���ڶ�������:�eʬu��61��n��)�2L�.�� ZQ�����B���B����iRw̚i�.S�T|p2N��f���(���	�sG���y�a�AZ�����j8��EG8x�O�g��w��D���M���G�����~���V�`�/���/�I����F������ ���M%���py�P�gp����4;=�x�:��N���*!�;ɋT�+���4/�U����b~e|���~8к$�;�r�����>:�~�Ȼ�����Rύ~���U"]��&f�9y �e��?Fr���3_7���x��6մ#x�o3�S�E�R�m�ws�_�(F��!�m��$�z!�-�w�۞g�h�֒F,�wY�5���jόe�nxE�i(�V�R|BeO'H9 I���:�9L1B���3��D�w��rgo�Q��Ɋ�׸��	x\��7�m�_�-�(Cj��T��׈�����XﮐXIȱ��������*���x��*6�3'���[$W�'�	�o�W;�i�Uz!Z�{��svc�p3�Be�vge'cd]P-py��"ă��,����z����
��v��V9n��<�3Z�=oV�D��~�V�����bh�~����d�4/��]�`�_t__KEV?��srP�3�$~N�ZK+ȵ/��v7��qN��v״�|��>52�]���Ϩ��k���Eߖ�Jl�9�DP��fjݑf�g�m��u?�S��$�gh��x�^�g��쫲A�.>t@%�,�l��V��Z��+<zY(xr�ϙ���
4����8���fi!v�����J��c���D�"��)��G��2Љ4֞m���dL$=3͓���pPK\�N��ڴ���c�Wŉr��W2�����~��*��s���Y�u-�&;"��u5f��]ܜ�n[1�!+j����w^�p&�����-��ff����؁�����a�:�g�L/1 �.fǶ���	�=��Q���_(:��Ɏ�R|�V�Xw-��[N���$j�Y�-��RB���]&����u$^��|������+iNU�vX�$گ��,m�W��Xg
#���J&�-y3�R^a#C��!�&'S�5�b� 2���0��&�h�O���?����r�U�p�����3Q6��0��ꈿ��8����O��\C��-�"I}�*_�h� �ʘ������IJ�mXw%��<�KAE{h�9�z���"�;o��ըZ�}��	Θk�M�=��� !)ϫ���T]���=S�I����>�y��ƌ��05�Z6��6�p���\E[���hǍ�����`5�������g2�;��v�%��X��dv0.%.�����l�qn��H��l�Oڠf�:9�2����8j��ʠ-cٞ̆Q�c\Z������ɣ�����M������S@3���V��yt�H�68�;*�����!a�%��>n�"��� �����#�c6������/�t�i����Bl��r�������{3�h�V�CL|��GVu����qз�c�4�2M�c��Q4p�/��&���@*�D?yڎ����:���K}Q�N��t��SP��/�T�>���R#*,���58��pJ�	7pf	��9���gԠ87[��`h�/�!�$ւ~�A��ө���� S�h�>��I���r��c�*�.�7�iM��.��ڍqp,m��X����"\:v^�EwH~k:ʦ�ƈ���p�y���`І�H��q?�ڷUm�ܢ��	�:�yq�!����`�9	��̞qp�p���a1��� x�g��-�MOo�V��4`x0��]ILm�����}�A_���\�Sm�G$@'O!�H�*�*��֗ߴ>�˟�|e��k��/P��r��;�=�ؼ7�{�P"j��8FY��A�U%�5��ق�&�ѽ������$F�4~�]��ߘP�h�O7
G��>��Աǡ?c������/YՑ)Q�?��U��*�ԋ�Ո�չ��ϥ�%�*�ۀ�)���u ��Ikp��\R��u^�a�ч^R@����9��W��o��;�#Bb�bz���`�\�Y�މ�g%�g �Y*�g㉻p��(�A��my<w��X�|�G��D�}}a4�&�<ct��kwI֔3}��������� Ť����<�������Ptt=UO��M��&�H�Z��ʔ?Ő:ܶx~H[�@t1��$
�m�|�([_I���H~���z�W��8�o��wp JXy�����<�����4sʼ���Bg؄X��$$��@r�Pv-N�����,[�fn�ގ�?=�S������	1h� b���##8�Ӏ7Bs����k`�M���J�l���4�x�1e���c�q&�W��ph�ݻ*�=�7�q��>��ѹ��4n���|��@��(���
�ϭ}��Y(����Aa�k�;�M����z�A& ��=�'��$LF��+/G ��s����e@//�?�R����*O=mt�yi�P�T��YxE��' �#���J�,�f9$V)9��[��}?~�?8%r50b>=}^*�c����q�Q���b���Knt*�P�r�K%B@�Ό� GyS����L�h�Kб�0���b�X|��h�-?bt�@�:��y!+N��3@�1C�5K*���,R"
���	a?�vѻ�hb�ᱭ9L��6K�f�bO�[�߳*b���j��?�L�1u
?�aْ���Xz`^h�e(츐�a@;�O��waƮXe�`N��X_ uf�oM��M%����y��/n�ɏ�1�B��O��������֮�R9��n����/q�]g1�ȥX
����P/#u�n5yI��~�7�־�q=JTS��:�Z�	|;�ϣ��?�g�?,�j�/�Ln�')W�]�:�"�r��R�P��/̝L'�[�v'>�V*���dh�~�����S<����x-��:����^3���=�AƣR6+f���Av{)���耴:�qy�B}�:
� ���c�<�:י)[wXZ���;���A`���(�$sՠ3(�&��K�Ϻ��r�ޑi/R��Y�� ���?t�^��pL�j��^�a�2v:s_m��0t`�:���K*P�!QG�Y��G��P[�/g�}�~���j�BN��7J��+�:n��`):uR�
�L����̙R)RF���Q��w3��b�z~Os��L���G��nxK*�IXȒ��X��2n���,8FUY/�=(��/3�0�c̑l ���LF��݄����X��u�=��>�g��Kbz��Tj�&`zG�X�w��D5��p6�qQ����BѠ-��e�k�aHwk�Eg=�["��d�Cg��w`��:X���!�1^�O�30i$6�"5�k�C��N0�e��o/���������܊�V�?��)���Y0�p��>D�9��s���ZF�ct�r���-\���L������@.(�&ύ\��u�Gj����T�Pq �E�SU&�Ւ�ư��#�"�-k��X�[����� �2�KL��͘�D��ka؇�^2r�Q�S�����kI�eV��o�)ʂ���'Ks�+6�	��P���ɏ�E��c���x�5x	Y�"�*�$������8Y��͑�ʱ?U�u�\���"�Ώ�_J�O�/��Ƕ�m�G�����2�����$�c}S�ҥ�q�Z���Y��J����Orw�S���(6��h���w@�A�{�=p�[�S�Y��|--���荤v'6!| ��L��:���&Xw���]������^�^�~y*W������A�c�������'�D|���P�C�h�yAlDe��~js7����(�����U`15K��@�s�RF/�4�l��Ƹ��AD�j[ߔ�� -�@"�:;MI�D.�������^s�:R=�`�����Ie |�h�|�����٤����8ElS[:O7�o��T�Ӻ�oxL�,Y➘U�n��/O$��+��	�)5�����$�P�:��c��D����¦���XSK�Qɦn�
wj��n���	T�KpXt+��ϙ.58,��:�uXV������K+�����V�5��p�ځ9B�U�bu�_���`2Zm����#&b����Ф:4Uِ�3�V����1YZl���[f�Ix�:[�"G��D_Y���z�c�3L��x���3W��g�	(L�y���6J����g ���l�!Mƒ�ܺ��n�:�y0t�aqd�����s5٬�A{B���l\���m=U�D��p��jxϦiSؓd�~�G	|\9`����CO���`�bZ�iR�����I�w�^�`@(��
�����_�ZS��?dK��9~���������י.�Xp^_g5K?�FJ^p�{SY�ȅ�&��Qd�g��1"06��#���0�0 _����&�0�޺��!^ޱ��ø�(+�k�k�x��17��"��^��mj��+�]����Ĵ���';x�ÿl-{ ��diϷq��t�kʮr�g;�27�X��pu'
��ST���ϻ��2R����?���B$3F9�[_�c]�,@�Y)�ԧqLS�;ku�S��'1�jk���nD����fk���U��w�G��5�[�-��G�
+�U��i[��{<n����'����N��Цu|AM��h�YS)>�O�Մ�x����fZ�e�NG�!r�Q�ĄK�7�,A�;@���o�<s����ț�*���u� 	�� �g-7��%\�4'�WF��R`�4�FCbw�Ŭ����׼�������&�f��/b-jq�t���d�O�v��[���#�8S�b*i5Q��b�.�yG!�����uv}��ڔ�8��}��#c~�1�pǟ�gΒ����c���^s�|�bo:�8�B�:mm�B�X ^4�:�_�-`��4�.$��$̬�N�֩����\�C����W���a&�Hu��㍧�=��%�E��1Hl��~�N"_�����Jy�H+�g闾�ԩ�,��'A6sm�o�����'��uS�_� �I���c�h����߁D+1�Y�뵄�MVnK���מ+��+��f�@(I*8��2�#�D��q�;+�>��z�`6�6�q�,f؀���W�jMM[q$sӉ4���X�bІ�pUT2�:�f�f�	����Fe��զ��Yt�hVTV��1x�c�@{�=N,���u�����lJi��X)de
�I7��A�p��_�>1���/6WV�XRg���¬�GB�8?5s~1�ASAj��38��y�G�ҡ-Wz�s�!u~Ӛ��֌�K���5�!y�k��U���������τ��}��W�L���y)@�dX�8�Ъ���QA�_%��yNG�x1���܌��#c �$���1ϔu,��Ϋ����ۓ>"�G�y�H=�e�e˄Z�{r��N{t�pY�b��#�d}�+lJē����@�C납��b�Wq��y����� y���e�t��A2�e�)�K+�ߔ4��`�^0�t�"%S,<�E�W�.I�|�T%�j�5��<�ƀ��U�kG�t�����~�e;�_��l\̫�z�۪R������V�[���1�#�?թ�qC�b�X᳥�E�~�DF�g5����c_�����}�F	^,cHF��D^��¿X�@*��:F|�[��p�*�4m��h�,Yf�c&aw}�4m�C��,�zY� ��hî�=�0����ZS�#x���b�~��E�4^ ��!n�ă��H3l�,��Zg�����lq{���i\n�2i�}��l�	�b�>T�c�f3I�ϔ=pܮ������j��������
h��h���4�#�Zߵ8��|4~e��rޗп�y�+v�|S�������j��/�3.�kNB���<N�c��W�����x���c!g�`ƶ���F�PT 3U�N<��T��(�o[��;O�����a4�㚈|7k�\�A�yyB���qg�rn�iu�{�
�$�V���6��j���յl��ɠ��[��`�ZT�D'jC�vg���*1*;��T�]%�P�F7��@oʎ�t��%a�?���	Pŭ���հM@�xZ�īS�Ie�����v�g��42E(;N��]���T_I�X��eF�q��[�6��ŘAʦ����J�3��E��s�ng� h.���z]����>�:Ge���z�w�ZB$^(ߺKt���?�EL�����)OW�{J�e��9��-w=	OͬCg��@��6������ �8��m���.�GWs�=�əm��t��:(�֝a��3��j�$[�_�[=���H�ѥP�T\j-/�y��]3�U12�m����:6?V�R�'��0�C��]�H�U-g��Gr<����<4��w.��h��o�œ����/�
���#j�U�\T��ɄXU�ڇ�uO�z!1���u��Q�
eyx�")�T����BhDW�"�=(F�4߲�i  2���%�
W!/s Wq�FT&�7 7�Q����p�)J�
U�޸�$�Ԫ+���sN�+Q|���!��~\��W����>`.�4l̗��m�fV��� �w�E�������p�ыM	�RN�~�*�NgI~9��b�W��:$}��4�/a������f�otKҮ]��v_��/��<�����>�.S9��:�dTl��9���jCi����~�Cޅ`��/3��������~V]���-&+�����̏�;mZ&rZ���1�˫3B��aYS�������v���~zBfO!_�:џ�iܣ!f|�vC�r�;m���"G���[|��IK���
s]��zQ�M�����z.���j!��o�Ii"���h� �,�-ؘ�rΟ��)s{��(J�ؾ�d�P����(cI��sR
�,��O�A;�����H+��zRԾ�O��A��B�~��v���G����/�7J��#n�HL����o��b�UՅ��όh�j%�1��m�$*�lL�'���K�p�vOZƚ�BS���ԝ(*��,�#�1���L)��/xr�ƾ�m1��Jr3���F���>� H4�_��bY��]�KҪi��> W�1?B;��$�0�r��>:T�����mzdއ����>�+-��tw�:E���b}��W��zP���H�(���Ͷ��,\46[��ٹצd`���jA��?G�CV-ՠ}w��������:��cCk��l�fu�[A���l�B6�L�߶M�ZIz�v���L�a�Y��E��=�i���6�Ƅi����M��>���i�o�\��_<s��۱����~��7��z*�p�}͹�\���C�)KfB�]y������oL�~�N2� ��d�n�9�a�]�&��bE�?MgC���"%٩�����·�r\B�x�DF,}a�I�ƀ�H�Q�����z[����"v��4<�YI�+^/�o�,sͿ&�exF�*�.	o����0�)��!tZ�~��_�mUF���gz���m��a�p�r��O��g�EM40(y�=�`P~ݨ��[��R��Xtmy��mD�Q�����(�U�Y"�gzdUߦ�z`������D0h�E��M��S��A�p�r�h���1vCb��Z����N3x	�ႰK��ot!�ѳ7����-���3A�qZ�m���u�7��P�ۋ�c�J>�Go���Ɏ��	D��[��ľ*��Me���o#�&���O�	-t�i��p���aѢ�.E}�ځ�c�A��W�h8����o���[:�뛧�B���ׁ��ɲ��a���w!�#X�$ݜl���J�-?1��6C���|J��\F�:<�0�6�MAJ��R����}t?Qb�@>/968�o�@�w�����roVT�ܞ�#��n��r�I%��]
�,jK��;�Búgb�euxP� � ���U��rx�y�ՙ��	��Hn���Mgs�.�XT=!F	��Y��(.��yc7���ʾ��_��� }���H���< F�3���f ��xB���qjaI��.Г�HR�.a���[3o������r���j(��uvC�'N%IM1������@y���&\{�搨�v���͎�q@�|X&M�Y	@S�A6��bD;m��fq7?\�����f�u~b��`w#T���}u�i�����:E�Ţ�Mq����e-�'RIi�O��03�O$�HA]�'��N�/L
������<�����ry `�j'���
ͼ���_5�!0��8:pN$����ĂZD�ә��[�e����
��!����o,��yXp�_��Ⴅ#!�O�<������&=�_�Lf��@�_� p98�H��*�ÈYixu�8���hu�$#���E�ggO���',��uL_���=�>G�U�,r�U�U�*��tL���x.��C���aP���� ��ZNl�JR��QR�Ӱ=R�Q��Z*/:c�5�ܔ�⣴S���[ 	��H�#h7��-�'�tF,���'/���/�ܞ�zl�v�8GP�.�я ��{�>F+y�����{@��wye���$ec�>��䞝��{i}�b�'��Pq�)��ؖA�!Tl��ֱt$����%6D��sr�S���`ӯ�49����g��˱��tcԇҝy#�]�����Ul5�K��H�~�A�۲�Z'ka����]����rs�<�dw=�yfx=|_�4����j�b#�NĴ����c����>�_��
�_kac�f��%�
l�|/0��Q��8��4i!XD���/�r��;��C΁X�c���ʘ�bf�XcgU~���� �C����g���+��������/���	�5|�S�|�r��@�}l��<���1�F��0!Rg��������v&�J�j������;q����(-0���1��푨��B�(���Jr9��^HVsJa4��ti���
W\�l�j�!kj��e�Y����ז�~X
�iJ�V��|�s����y{R$�"���(��;�B�`���l�k�"N�8�,Y�N&����T.0=R!�p6�&�ʥUo��XjӁ��*�n��NM4��$����E=���l�&E�ĵ�d��?���zD�}�n��m���.4 ���[a},�~�<b��e�nG���0�ڟ�M�\s.����[��K�641?׻�^���}J�~;H�'�S�$�qƋ_ؤ����Hڶ!-Z�0)��_�2ٿ2+�����fR�ߗ�i`�x��#X-���aȜmF3��Q�#|')���׆a��D
�l�p���Y��d.�e�9��k�ݾp��5�A��MMҏ�@87�k��q[�Λ$`l^��_����:YA��	�ĩ����e�)\��� �Ͻ.�ሔ:��~n;��%�Π��&��W�i��N���9+�w������4$b�y��N���z� �4H]3���>)�1�K������mXJ߹��s՘�L���[6��'���Bﶂ*=�:���i���L�$r�@�>k*�` �(�U����W�%�8����JG���0���>��O<���b>M@���Die$
.�ɁC���V˃~,�^Z,*�s`c'�R��R����sr���&���}�f���
L�L	hC��}��e2�s8�w΁�ZT�;I֌S*y�}	A \@���76�M�~��\�k/�rNJ �\;o+�>h�xrD��r���v�j31�j�Ֆ#�@X�Z�-ȷը���o�}e�_���Y�Z���1����ٯ����&�\��-��Tw �u(�'�Ⱥ|�=��"�}���M���t��Z���D�u�:��>�7����\�;l/6��T�sk�X:��z�B�ǉ�f^Mi�wV��Gl���(x`�_�F�D��aJ�Y$�������m�~UhI�����ڒxqm�����-#�OF`f���X�Y��{�^�Z��V�1��?�W�������sթdS�����0�V�w	EG+^���x�踚�f�\�x�Xa'��]�}J���e%��~bq�O%�W�=]�����Yc�H�?= ��KZ]�[�n�������a������2A*Y�+&,�Q�Z�_ ����4�ظ��չ^Lٰ�C�!��pm$/ʴ%��۱�n5����,qHasz�Y�g}�h�a��.�nS���R�G�wf���E�y��(���R��E�@Lc�xv^8I-Va�a�����TM�h$+"1wC�3�o��!���Zc�G퉍=��Ԩ	�WpF��q�Ë�w�uJ�����X�FzY�wG�#�o�������i�t����� �f���`\ꅢ"�y���S*��2�[d�.�k��2�
�����q������0��b.�%�Sd> ���&ނ��������L¾����}T�݆.#s8�Rl��1,�V�����r��[����&�E�쒴Fp��c�Io�_�����)|F�s�B���6nF��g/s:ڭ-�}zA�f��1�H���ـ�9�~o�3��>!�L�S[�L��5V,���`��d��s��ɲRm��J\��D�����3O����ɮN�3q21�2DNH�l�,y.�ױ��!��������:�F������E*Am$v�2u.�� �>N���y&`���!]Dŗ��bV_�|X2ӸL�mk7[#�f]t��Qj4�-=����Laӹ���A��(�<�/1�:8e���\0,f��By��YQ�s�SѢ�R�?�A�B���~=JȺ��+Z��1�6�C�J8+�9�}�Qs��޿wƱGֻ����|r���׆i|�)  �d��ޥ���	�d�ŭEb2B�/Q���������Xv ~�+����
�]-�F���C��tO�"/��ic3�>O0ALã3v9o�>972�ɳ�Vf;�b�v�Bݏ*�Ꚃ����W漹y2�����8���<�^f0�E��{P= "MB?(�S��h/�����S����aJ3��=��kN��:%���S&(P,�+��[[�	/N�}��z���V��En�?�|L�U��l
t�l��� �%y^��G���Z��P�x �q/�N}ʃ���^�tW��j�i�'���ﺎȬCɚ�l��r�uX	6��.����V��4�+Y�mQ�)���7=�~yH!cY/�Ɣ�49A���a=�PG����L%+�}r|"���~'�<�
B}0ގaJ��w�hJRs2�޴YRt���c�|3��̆�{A,Ƶ}[���^��>A!ѻ�ov��wX��?�� P���V;� Q�\��q`Y��Zs��O�f�lo��{�LŊ��f�%oP���Aժ9��7�����s���񊷦���r�?���v멒��v*�]@ Ww� ߶�`�$�B͠���5PC+���Lf)i�X"Y�O��XQ���kO�a�4Y�?�1�q��d���l��U�
�������y�`w��	�����Ld��_�]�uK �e�cH4�>���o��|��i���	"nt��� I���O>�J�h��������,D���V(ȩ��cl��.�+�Ŵ}�Z������ݳ��
0y��BS����)F�v���F��ϊZY�I��F"ǅ��F`�Zݱ�DZc^����f;Uv��FD��B�a|�VDu�)�~H�Q���kS*�Ă��{�Ij�ou���5�+��`_����Q��z�f�}G(8��F��3��"3����]S�?��+<]c=�G�C!'���)�<˷t:kVa��ܳ�Z������	�� a���(fD1[F�rA?x�#a�u�N���^���Z�]�ّdOB
x���5Qw;�UM%^��^��⏵)eW�cA�������Q�՗](tt��¤�%K�Čk���	S��U֮�ob���y'5E�T�����M��(G_��p1������s-�3߈N�\{9� � uR0���K�����k�I7eOJ�\�Y�y�B�,#:��	���0���Y��S�/�ı�۞�~�~�=�Ec���sfs.���ZUT�15�;֕��d���5��*\E8'��t��fWpH��eX7Ո	���r0j���sT��YT���5�LCSR	���F�ۮ��J��˔���^)�W�2��!i�<R�2e���F�h��Sn�7�0S��X9ǯ4?���P4)Ù�Ba��Y�5��o>H��2�.�n�U������d�A� �0骓��O�i}�?�)[�k�䣶�ɼ��Kd�A=R�WK����H�^�-2��G6��J@N7�^�����Gp�WZ�D*I�:�E�u�E���=�\k��g{�S������]�I��+m(��"���|�4�,1U�Sؓ�D��1U5�r4�x�sYy������VĊ�BID2.�m������}vx���q�/�*�������Z{����
���T�J���}�2�Y�����-��W���}̩���o�s��S<�$�0ZC�q}�����u��\���٢���J�a�\�
��W_W�_�����Q--�?�Y�6KҤ��<uK0C;�0N�,�|�*�z�pT? �G/�������2	둱q��k��8(�G.�y�Y?��
����e��E\
�IY9�u3�6�"��^��n+�"��a����9��o�SM̅�t� ��׌Z�`0qY�3+�h��8�4���C������%&y�'#*!(���剀)��|��SV��څ����}�o�5��!�@�#���NxA&�������K�4p��,V';c:w��qQȶqn�Z��$��-����*l��9�?�k�d[t�<(�x�/�v�!�J0cKzn=�K�[�\��a�|��Q����HP��>]�`�ct퍘��K#�x	W3����Nfl�d��
����8u�]�o�����i��&����������˗��[����$a�+��m��m��F�UȩJC��l��E%�V��4'�a���J>� ] F�kr!��*�&��~$iϊ�M?K�#���n�s	����\��n��yK�-A�x
�Ò|���Oq�5�{L6~��LAIzㄙ�H����V���a;9����W�!S�����0Ѭ�!�|Ԅ,+�S+���݄ e傫 ��:Ɇ�A(�����yF�re�m�B��c<ɛ�m��ƶ�k%4�P���]_�Y?�(V�DW�zg��	�#2�˹����V1����W'7^%)N,���Bw�1,�l���|,��-�����G:�4�����t�nV� �G�Nup��K�-<x�v�}z��<�<9�������a���h�t���Yr��VRT�`� �3�
CE��)�J�i��#;�� �N{s���J~{ ڭm�D�jt{��y{LaW`76H�m!�\�Ɣ��=��"xmF�5]D<��W)<���:-���͆�}`�K\�
��:�ު��(ϓ��;�F���O
T#��}>;� �%�g)n�堒dP��%[h���E��]N���k�4L�#t|��	�A9F��j��@F�p�F�� ��2�cV w��@n/�E�ݑsN���x�?{��������,��2�9\>Š9�!P��m��K�:����W1,�c�R�[:>�CU-��P��M@7�Z���=J)2���Pg��0IM�{���TBoaY���q��=���8A�'��y�x� �[¶��(f�� �|�����J�����M��t��\��齿����oQۈ�֋� �s3�����d�ږRjb��Ws��`���[�e�E�cI	A��D>�n�_Ij���]vK��� �ی�{��|V?�$R �s�����e70c��������������0Ȟ�(W7���R����RI�=0���5��8��ٙ1cڔ��v��t���E{@�s.�����Q��}���-�f$��>%���q��Uf�q�wλ=�e��ꃊOI��91�t�;��e��<��{Nt��ߙ�t����(ө��yMn�?�����$����bE$��8�*���cQ�<|f�96,�C,J`O��QH��[s���B�,���_P�J�w�&���L��f���u��U^��CZL�Dg�W��ZZ�ؕ��PM��"�!o��G\�9���(��팮	w��5����է��rq�Kv۾�Y���;��~�~�C}Ť�q[��s���Jy_��� ��\̒4��'����)4��v+�(���|O���
��r�Q"
�L@���/�F, ]5��Gf��Ԇ�W|ѯ�vb�A��Q���a�Iͱz
t�I�0��[�z!��
���D��D�)��t��!����(h���JOtf���LE^�*��'ށ������)�������#ܞ����~# ?�6�+	��]�?!�$��\��\6/]�Ħl7�8��v��D*ery�^p_�z�@j�Ws��vM�=���&h����.@�������%��}+G�'�JO���)��M6a��h�+O��Ŕy(�7Ed�2X�O�I�C��~�?��+��- �o��"[0�@��o�c�0m�6|�E��ư�=y!q;	�L`�7?#�"_W80WQ����ʿ�8��]=��](�2�Z|���Ju�*͉@�p���mՔ�-�ʴ�7Q__�"���Ò�X6?k�ҭ/����0��S��i\-�"|�k���?S�y�*�K�q�O�W[3�~+vR� }��E}J�c�i��t��}�c�x�غa����:�����tg��λs|!a�y����o��k�<�+�#}<G�Ɵ��%�Rk�{��06f�*�m1�ÛkK2�����:8N�:Bⓢɴu3n����	�9E�J�K�si/b�������v[��t��K� L7�q>���Z�'8C�6Y���zXH�%�\Q�3��!ڍq�OԲ4�{s^��u��~��rN��S�}�&x�R.X�1�laJ�j�-!d���{<�<0�8���7�S��ڂ����A�D�27b�2��lu�;���f[q8�y�WIJD�n2"�1&��=
�#���|:���	�m+>��bkWZ����)��`�|g����^��N���Fg���"�C�2�����E/�:��j�).�(�`��|s_^��B'B.��mJ�� �xmaP�zH�=>������-�̈́���l���X��F��A�fȦXk_��d�r�y��0���\u�غ�7�֊��X:�o�\t���Ҹ׌�C����$(;?���~_I1�p�%t�[N�����%�o�o^�4.���$ifXZT��L��F�(��ts�i ��Ꚑodd ��� ��Ph����s�!��!�_�E�؆��whw�s����n��
V��~R9C���jB�ghO��wh�N��IPVG���v�NIU��ר���#[��l���4x]%z��i<j�ѩ�خ��v4�
-�j�D��� �~���k����"�����~�zbv�?N�9O�����}Rr�xx��џ�2 ��ܞ��rk�`�ʀP�]0�̠����Y�f,^�݉��|*w�{*�9���T�ß'�������_ڔ����MܦΖ��\&�B|���t��^�[�*W�O�����ԗ)�e��o��.Y��+�$~A�(�-C!����=��3��[b��B�~�,��C�ZG1���w�F��N���觤/��_u�!���E[
��I�7�K'1�mٚBy&C������B�9�Q4j�ʇ��+��<�&z�]i��ԾEKLj#�N��U�Fs��z��dczQ���b�=�q�]��?���7n 3���ܼύ:���ͭ��!R��i�hv���4A��ɨsգ�9� ��.ˣU�Do��e��HRn�:*���F��� �xl�M���]�@��x�Y�Q��$�:��jM���y�"�S[�_��iR�� BLw�����ǒ����`��ud`���.�l��1y�n��)��Pj8D\���s�������	��R��4�I?�VFq �W���D>� 7LA�d�!����ı�F� ���lY�S�7�υ@h��N�~����n嘖t[ >�J�Y�q�;��(�3��/@��~�OQ������x��]h��ᏻ��r��e��mĔ@�ӦsA�g2F��8"]HEh�Ȯ�mʟ�I�I
��� �ǚ8�.��XzX�q���]9��2n�5��jQ۳�?P�(Q�u�#�nL1�_��t��>��>��W�Ш�;쥾��8��b�:��s5\*���_���Hi8QS�Nj0e��U��GE������4;�QSt����M3��s6��Q�B���jqf�m+��A�8��e�k�i�n�^�c���o��9���._H��4��ӣm�JT���"d��=�Wfn1�D��(
��4R����&
w�)ɹJ������o���C��[-�_S�����j�pe>_1����!�5Hg�'3�7.��E���^��ށJ����L�3T7��u�����jn~�S0���4�E`:���?���%*}D"�iU���P��<;�oU�Q�d�����?�{<�C�Zw�����S��J�o�f�i+whyy}���'c2; 2��U��$�2y��`5j{.3B'XƸ�cSAhR�	.(��ہEs����C�:K���m�Ek����� �&	Ҟ5��?�Z�z�(� ƿ�m�H�bn���y:42:bpB*��`�b4�����,�H�S�[	���9[8,�7\��{��d.�ĺs�ߞݫ�Q���{+v�mAvb�ص\����%$)���N��$��� 6w��4���l��bZ%���8��	�	`L�m�e(!l���PF�&�=�װ�>?"~ �jג��K�8iZDKe9����[�0]]޳�p-��.*���]��tQ��n��5���'u��>�=UİW̬���t��X��j����8Z���c���%�@��.���d�?�D�ٙ��.���$�qn=�Q��p�Nv\K��S
�����f���4fC��%�\���$d��!���S#:����1�Nj����܈��������jd;�N��I�Q�1*a��+\���$htL��m؍�˺pX�qτ�~cʁ8���(�FC6��q�����+?V�o���C��5��F0��;D�}��m>p�\bn��,��m$��L��g���:����A�L�ηU�S!�HI~����R�E�P���bCp�[?�`�-d��R�5� 6��8\�7�v��V�o*s��sc�|�v���Z0^�s�<�RLP�_����իJ��F��
hk�vn��͍�Ur~�G[�@<�o,���S���j��&���n/k�&����<�:���t���`��%��A�I�0\��r��AӬ[L�����1-��Y����܀+��I�]�yCz`w �V���>^7����.�����do�Y�r��~z�YRB#�Wu��Z�!U1�a�@��dRFn��$?���",�1(�`%k&}L%�� �mQ��C7c5Y&�1���)�hf��<⹰��6U��f���5�"G�V+qYK��]S�q�Ei�--x�y*~�-`�=r��F ə}I����"����N��|]�iC��@��0���>�m_�U�.�@D�o�3��j�ՠ�A�������ʿb��6�����as����7���P>���T��Ͷ�5֍E����V�����;��. ������<tx汕����s���A�訚�~(Nc�o�U�٭�A��R��-� �02���C=#`��z�vC~"�U�_��'��=��Ԙ�L�+V
B���˔hW��H#�����L�����(�V�$F+�g�����Ҡ7-%�!�����,{�x��-�G�?�&X��t���.��w0'�!��&�������F�Tm��E�K�A�a�p�(�p%'�}�~[�B�Jq���#8۴P��V�p31��P{������hOK:�PQT˿cC�5V��.�M/����K��@΄, $�:j�R�n�/� �7{��V$r�MAu�2��S�GNr+;�)Iu_W-G�r� �-�i���s�j֟l�м����4zd��(�������𳐗��0����@����,�;�e�� > �����&~�9���>�K����HB������Rth��&ZFN=��k�gҠ��k��L~B`qB;W��,��*�$Ȋ�ґE�{�R�r����L�E@����V�
wai���-3��L+�]�]T�)[��Y���iP�u�ۉ(�12�� �`��LL�6�Fx��u��ÑD�׿g�����b�p�@$6��*�#��2Yk���?�Og�)�B�;b�K��e�Ҥ�D����4��D�)���g�nCv20�<EZ���XDE��B2 {�fCG<R�B���B�����q�W��3�
���b8����R�W81EK[��(x����q��*8�d�6�xs��?j���-)��^�j"�>�#��~q��Z��̘2�\X�q����FL�6��p4�l���B
�Mn�\F�]��}��'��f��|�����E������OA
>1�Dl�R�ol$XY��(�R���m��c��qZ�~�S�;�X�ׇ�����OMT���\���T�t�󛮧���<aY�Sc�������;}sG�*�o�\��Z=F7M{�;Z �w7��ئ��/����N�7}�7��(��OrDi��@�|�=���,<m��`2RI�F��3�������s[U�N��������WH��	�U�b��4����b�SnuS�U9g5����V�гr�oª�E8	$�8	����~�Wh�B�ԥ/�F���O�+@�C���%86�j�X*�nTc���P�t�9/��Y
z��o��3�qk*`�����8d�c6&�0�c?�S��-]�#�i^��M��Qog�X�R�� �a&TnOc���iT��4���Hۉ����$�On��'��r�h=�x���}O��֟T�����1K��|��I�� ���[�ۀ��6ޖM:rK������o��W�z*���VE�G�?�K��Y�*��{���{^��1�Hr�EG�ҵHj��J�>�19�ސ���?�
�J{�DV�����o�<ny�K
&z�䜖GhG}���^�#"ʔ��wԪ+�#�;G8 eҾ��A+����AA#�ܟ�G{�)��C_��V�����͏�|������#W�diF��B�!��_�N�x�� �k��K#c_�s�0{��C�e����H�D6)8T	Kg��H��g�o�u��
�$��I��m5x�h�i�[��K�K���],Q�M�u��q�qd��+�>��]�H��jؑk�G�Ƙ��Z<�ܗD�=��V=��{�fe
1���1�(�� ��].�4��P	�!��Û�$�VvtZCMw0��!�2Z���y�٧�l�^�k�:��T�d=�K�rq �����T48���u@}Sy�Gŷq$`�h��
9P�v�٘ĸ�>�
�^SwW��j��W-Jb0(5���I䐚A�-3����l��ñ����Եۀ�u�y�u?��lIC*c0���4�����y���m����/�j��JVp�j>����|�&��]�ג��Ֆr��cB��C�N�ڍ�K�?�vl�4�S���f~i���t,����E��f�XstY"g*>"D��e�M
h�΅�D5X��Mf���g�+���,��n�%��5���C�ѭR)��X��P�0�Y�k����JP�XUk���W�q�(�~�����m6�ݨ�ن��%Ý���RD2�<NQ<58�������g9q.G����kL���(�5��Y)\vm�Ӻ~8���ڟ�/!��ꃬכ͵�Q!y`K�_��!���l�5����j����t�%z_�)F��΄\/Il�v<w&�ϋ���B6!�u	ߵ|�=4�2��WlW)IE��t+ 5� ���,�ʀ�.��wo\�ݪ����7���5��"�λ��O�\Qg{��k�Rh�7������3v�)j�?���{sY&k���!�z�/H���Č�;��;����#}�-D;W�П���.\��lʧ�e�nT��P�IV'J���Ƚ�4����������� ƕ����t�K.BO�������H[;z��ˠ�,kO�p'˔�0��-�*L�����G���6�ز�>ד庠�ǩ�ѩof�ɫ��;W��gΑ:j��-X��K�d�,i2'����z�i�٫h���l��K��o4�z��K�)���]u��X�R͆�X���5(5h�`E5�ӛ�k�o^)g��ES��.@d �h���Ǳ֪���bX���3'��/���Hi�9K
��lU�FH:�ّo�U{N3E�W�
:�^��j���Z0Yj���@-���gV�1�?����S��xNye��\ܬ�IL�rh��FԐ�JL��9�E�E��p�N��=z�=��ʇ�V�cmz%��9$s0����i"ܣ�y!(�3��Aߧ�VF(F�H�Nr���~񔃝�d�O��@̎���Gs����A��0f��`!�&���ޘ����	��E��� �;�.��'1�4ې�ά� W
l[�D�M�5�2GH;uE�(d�N((ʁݯU,�Jʶ�l(�
&����9�D�m.���+�t
��u�b��
7�_v�-��}*d�Ih�{%np��o�q}�1���0x��<@u�F�E��y\9�`\�
�yV�u�i��W����8U���\����%�g��"^�Me��rl�ŔM\&Kզ�0�-�o�x��,�̉u'��^�\���_��=��!���\]4:�,4G�^9�g�r|9~RE���eڸ�|�G�,�Vy.Z��7KW��3A�O!ϰ���W��{���(�� ��U������±���3��y'��Ak���ӤTy"�i�=MLf������,�]MP����-;/vB�-e0��b-m����P��+���6�)�	+	�u��5��6��=�����;�Ob����V�?�����Fp��N��Gk�kŜmUƉJ\D�_����\�cOU����'T�a0��y��ԫ}��P1nv�!92��� ��ە��uk]��
b�ɖ�A$O��n�����%�?x5����Ϭ�c��-T7yq�w$��4����u59)�Vq��4P��;� ����gu�M�f��W��Md�V�Eg�Y+��0s��i�M�F���Ve�g���)��6�:�C�?ά�xF��~���������5�` :<��Ь�!�AU��;��6oo�S&%t���%
iQ����S�A��������(�{ɓ���טs�c������3�1������,�Zi�5��s��Ij-$�<�pb�y�Ȉ�����9% �f��1'VOiN*;�@��#}1r���[�Fx:�#Kk�f�{v�UU+�I4����J��F|ۛ[���͡H������O�p����D���m��d�	 ��UK����^(I쪁�ian�b�Ϯ�
�(����i�gD6v@�^]���/�z��J0�a#�d�g`�������S@i�O�gRa�G8֍��<n��Z�Y}�,��&7k� mOk�ٔA�y�)K�cn?�Zs��R��5�x�%Xf#|�1D+a�� `	�9�H�kkc5U�L�+r�~��P��O$�vkh܅O���
�-�O!%�CP=Sd�O��E:���S�c��"V�f����$Dq��m�S!1�6��I. � ��!��!Sk�4�x�����ˉKs��Up�G�N�,��$�¾	h&O���\�v���2 ~���4g����pT�U�i�����st/l��������4��r����/.dA�G�� H"=?�Wz���&wGǨб�����_�����O$z\
�Zks��_5�Wg	r`�����ޠ><\}m��pv�|!f���Bu~���p�~�]�c��p0	�t5�p?�쒲�ش"�q4B�i"�8���9�	@�S���}v޶}ނ�ގjA�B��X����r
"�P㰧����m��4��NZ�����RS[�a�z�yT§	;�Р��*�iL�����O(<Х��M�쉁= ��TA���@n��i�=J�g
����;�$.�L�,�;�2��N�?��p�ե�!��@7��H_(1,��}���]�� ���u �����c�A/%�
��������H3�K��U���x�nu��}���UivpWN<�.�J�;�U?�01/�C���B'�Cu7]�m��
<2�%��-�Q�a�!�kqj]�F���a�e\�<��ohu�%���� ݄����fH��~n]E�����o��eM
/�G�̟�e������5���{�^�Mz�T`�#�f�Z�c��A�M��_d����\!���L�E�����I�)q' ��q:�o�ؖ���k�<ΓZ��q	V���H�ĳ�}pq
�	�B�hsHs�D,  �մk��n�D|�P�^����GA���
��
��W��嗮��V�Xy��jM��;x��W�Ȉ�!`	��|��7dҙ��2�X�@�ݔ�r��MK:�����jH�]3�6�����+^���R<�YԲ�"��Pò�vFL=� "=��?uK߮�Z��!�qi�f��6��{&�ǯe�*4E�L��sB�ɓ�W	!�����^�ۅPd3lxڌ�5@*|�����3�lI����?�ő7�Y�[{������n��==�ҡ>[�)��Z��i���U^��d�ý�j����ao-$�ֈC���y1'�~����A�K򟔉�G�����*;��=����!L�u���6}���IM �\�w�ȔݓG	G���K�b}��^�8H���7u2�|���C4�8�w��Y31B�.@�A��0���%�+E$v@��4��1F,*�t��p�1o��Ӓ6!W��Ğ� �`�P��ٝY����r�<x��/�C�y�MY�ۇ�SP39�
�v�u���i(���5d���pe,���+�<�TK����M7�ȕD܊U.�Z P��R����=��e)��
���i�.��":�����B(���d��+B�,7����=��扜`���aA����UA���f�v�Eb؟F��$#݊R;���6?�E|-J�W�H��%�*M�Y��������K�[A�Lˑ3J�.�|edR��k�,�{Vk9C)�q�T�!����\O$*!{���h�{��8����Ya�,]3YI�3�d���<�b&�P?W\r{֨����;r.U�dĨ���ЊS�|zJ�7يHôr���=Gw����%h��>�����gٹ�q�����sb������q0������c��}��c��'�"ؓz�K0_M��ܹ�&�j� �"��+�N�J߂�A���3FCe�[J�͠��y:.��$�i���߱L��O��U��D[B��c���<	C	�J�_]U	b+{il�adA�5��|sGX�[lӤ��pkce���C�8&���C�r~
�<�_p[��Qh��I�̨x��!��@�L��� �>�|����de1n�F��Km�H���
�x+K��j	�ƀS���wM���^��3�@|6P5�=p7�_��ﯹ9hB`{"^�P5ۺ9T���ܘ�\���
�L�iK�k)T�{/I/�x!|=�>Ъ,ږ�0T*M��d[�ד�b��������)Q?{��ǔ<_��,4����:I���Z��:��p�zX&�����5�a���|cd����]2��V���Q�\W�N)��i�m-�}�m��L��"��^2u������8��w*}��D�N�!��q�q�ǩ�_�ٓ�/
��؞؜�4�7
���3��V���&Etl���[�����1F �k�"qQ�,�	��G��|�E�
�Gh������,A�zd�2���4�D���.�艚yb��S�葸���d���!�0���������-��/�xI=��:*�pJ�Dbw��H�M�݇GqjS�B����B�}l�A�?aG�f�ȕ�*_,�սQϜ��x�B�D�S��ԝ��FP�ghz�lp��8��[3In��>#Bf��XU��e�v�&��>���(+�#;��y�C��x�=k�I�������M|��+��$}~8ap%ö�?�x+���f�ܝW�}iQ:'��f{��-C'��э'��W�ڊ���
-]	��(e�8��QB0>��bM��|=��f��iO*y��C�EIt%1��Z4&�����]���1��a�F�L��UN��<�<A��׽�]�D��o���]�!v��̎YD����z3�
�z�[���|՚�b�Ũ�(��NX������VGEUD������2���՗�����q�6��m��v,hP��KCrA�Y��x`�U�I@�;m��1�`��j17ԩ�$7��|Q	8-��r���p��A��Q����i|#h�b�e��	�5�����vFHj��MJ��eT�іP�'��&z$�,(���-N�~�k<�ȗp��g�	v=>�����.�����S �G`uh��?G[�q�W���1�5���VD͵�!R�ʳ��\��I�ԭ�l����d:�g|QmRi-��Ɂa��Ďtw�����h��A@���ށ�&�ʯ��f�E�~6�]�4$��y���kl;]ttA��.wu��1��l�t����p�d�6����w�j����y	��Ef"*���^-):y�W<�~�9���R�}��'�\58.#���-6����խCYaH�X�\�M�?��yȲ����Ek�{�	��L�#��{ V���r=�5
�ѽS�����QnN�b,���L6��0dL��I�4�|�6�H3/b�����.�1�ÿ�2i����/1	Z�20�Wy�$�$���5�>��&��cH�]�?�VJŽp|3a"20���W1J�����'� 4�� �6�Ћ������y�-a@ӏeO ^y���Iiȅ���;@w꧵���Khټ�]=S�el���a�ݨ�~~[�=��;_KF��)��0�[�_jT�k��'����-�����\�~Pu;j�⮖,�k(��"h���!x0x�!fm<��	͛���N�8�]ס��_F�;ù1�%%X�as^k��{���聍�(�G�_U�'˷ Jv�#�t�8����D`�nH'���e�Cγ� m7��b��|:�5�j�����θB��*}�.�-mZ����d����Ʀ ���,CK��_U_�M�{�N�N�d�<���EeWn�� M>A�+�n��c;d���#��5�~��N������r�E6�kh�a}��X�0؃a*Z�[��N%�/��j��7��Sr2��D�7�����J��8/��1�`@3�@~�jz���F��e��QT,0�9
��ua�Bȱ(��������Bw�Ȁw)U_Р���vջr����Z��HH��G�K�\�-�[�y�rU��1ȼs�*	k!�!�|͂s�f/���7#n��cTp����'S�i�ݕ)}����Zp�3���6�{2M���AZ��-�X!P��qr�K��A\X�'k��ڷ��=�	y��2��x�-ۋ;�X�Ry�D���qg3��ZV�PrC1��-�+ W��)�X�����:&K%�K��G��7A��	�!�.�j���,	�nHnnP�)NWsB��Z�m7f@+�i�u�����M�v�Fm\4�$h�P��f�,��-�����?���t��9�G;�F�����luŭr�R��BX�Ԫ"MK7m`OV2�j^6���e>�\�)�n����K$��k�SS��_p��������?����&U�����w�ӣ�IAE�8��t,�� �t�}J��WQp�_OX�Z#���:JF:�xX�FP��lL���\��5ОSb��C��O�|�d�^'=>���<��~Dn�D���}�ɵ���)�`FB�-�4�X(�YFfE���[��;Hz�*W2`q����X#@���}��虁hԵ/�5��y�pV�x���,&藦��Z�Tf�D�q>wL�m�k��N�/��A�Vh��sp���P��K��<%��Ҷ�E��=�@��8���������wN�y�ѿe�z?�ގ����4����X%�B�i�Y��i�!@:��&�Q&��MPa�Ic_k��)9k���W�%�~d9��,5�} oD��ʦ�ť�9�~�/����6��� |�HI��X���8���S���@S������N��e�H�30�/���M0���ә,�����h}�E��M��������;q���ï���Q��{0�G� �����{ȩ� ��1�^�-;�/�M"ɡ]�3��AF�ĩ�*�%��J�ٲ��j�������s��T�'W"�}��X�z��t2W7���ʥ:������݀2�[�*-�v��'���9l���A�8z�{�L3���/
���$������ �܀� ��H��%�a����{l-g.������ϴ��7-�[��,�f�m[�*��G�����:��]ʤD��mp���4TY�����I'鏐� ���9׼�?
UZY΂�J����[�����9�̄Q?���˚����wa�}�d��2K:�W,&�����M��]�(̇k������R����ߡ�X�D0D��f
&P�{~��I�P�mR~&+��H���V�٪KT����0�􎤷����Ɂ����|{g���@�p�C�� W��� ӗ#�W���<�L���_j����<�ĺ��z��̪)�H�t�5!-��uW�� ���Y��Y����;�rE�㱶|��4�,;j1
Vп :�y' �O�n��ju�ʵ��+����Y�<[+�r���X
�$x��)B����^�_J�����>��pߐ'�'��]B7Nu��y<���x��)b���Ї��G˂�ũsaUKt6�{�@��1�4_>Ȉ�Z!�`x\NzG$��u�d�v����������F��xf�N�8d�e���L�-�Oaf����U�(����4'z���E�g�H}_$����]��o��p�L�-��X���F��|������>�&��$����q��.���f?�/�[XA���i�푶E̾'k��> �by����d�����l/xεE(���B��.r'�@�lܰ"A����2�y�<䡦�	�J��޾��-���莎8H�r�$��K2��-�+0����6���y 3ς��H�mN�`�� ����^���%�Th�pǪw�I$9,vz
G*�IjWj�Mn9���� �����z޲�=?~vPb�(��]���ԛz���8�"!��[����|<�}ښ���B�I.Q�3��g�1�5�䂇�5�ڿ��S�����*���8�EN�y�q�SN�H��Lu}���l��g��0{���;�
+o:>S󋃛�t��C��'[��Zre��!}���-�z��4��&�m��4�׆��Q�	�˭d��c7� �i_5f�b�
>�m/���`� "���#z�$��� ���u�E�':�ɾ��o�\Z�uZ�;�)���E�a����m����A��M���Й4$��VFf��q�E�u�(��[K��e�YGAWY|H�GG��mS�r��R���H�9���=PS��Ɯ� 5�r������{�"W�_�eg5��Ƕn{���A.#[�+cC/�ssJ �2,y���!4�{���"��0�!�<�թ˺$�1�Z>Vq�}#q[��9����81�=��45@�#�bY(�e0Dn�����p�T{�[ϰa�Ag���%p-���Bb�:nH�y���+MdI���-7fGc��/����1j>�L
�?�~{3-��F���:��K޼����lk
��	k�k�L�d�
�?��%xNYp����fkӜ��;J(�a��ꀼ��ڟfV[���|��o�?ƒ�4���Ə\��ob

vh8���N��z�3\<i�޴
���E��Hu�Jd�[):l��h�	,��_� J�Fi�b7� jB�4��Ig �vz�ы7��"娱�\��͒�V���"��?���â[�9�ƒ[G��qzl�
Q >yÀ?�����. Qu�D�L\q��(
gv���<�}�OT����DDU:���R�?�V�$�f���P3�uTM �[H��9���{�?Kp�j�/Usj�6�C5ܨ���ҷ����J�H(ӄ;b�Moqi�p�dtmA��u�q����8Ɓ�|�����{�8�x&�M�!ɖ�B"����uEd�L��4IQ[���+Z����N~���ʨI@$���J�ط-�-�Z���A����ܼ&ٚB�����ޮrȏ�Ԋw�}f4l�t$7A(Ck���(�)*�����'�MÇ\f�3&j�.���_X�ɛC5@�HV��'��E��t*`�t�l\���Tf�E��g�w�W6���s62U*25�[�B���4d�z���g�[�D^ڷ�1�^v~u��bb��P#몛�> >o_��'6���쭠��j��WI�E}�U��1mn(GW���>e6���f~�Z��~�-jNĎ�Fs6����۲��.V`|�;zcҧ�r�f��Q%36��x�N�ʑ�88�=�o�|�i��h4�U����F3�#!7I��=?�������7��B*�:8���V��m��o������[B��}�!7W�)�̀���R
`�v���Iz6������[쵿�'DK�j�kނ�߄i�����Exu�%��Yj㚦x'咖�� �1vu����^���հ<k�o�5H�&P7���FUpC}&m�d�GT��"A=�o��W�nE�zXG�AT��_�~����z��݃B���H����%H�i��{>�+:󦚺b���@��h���,�7�h�F�W���	 ���󢂺���\��>��_��P�yr4�
8�c{��L�8�#� 񍓲�OD��/����&�،m����z���Ҫ�W��B����Ix�F(i��.��Os
+�F��w,m�.�o?m�v��.qVxq��uet��� O&��(�_�Ѧj������4]#�	g�DH�l)GY ��>�:n>����	a�)w�q\?EF/-���#g��S�䲐T^7!dJ0.F�	�|=\��\�:����Y���K�^(Â8�`J�<X�N��>G��Y�G%��ipq�}���vɽ�l���1�[
(�gܢHyyGH������;AYj/kw�_c!���g�[B�<8��$��E�r���bH��o���� ��¿�󫜮�����u�7����[T������}��x��6��p[���\�]P�3Q,���X�dl���y����Ĝ����:?��\�{����c6CcB�n?�d�h�}��8���ǅ#��S��
ĔL�5x�?��e���v�a,��n� <K�D��o��߭����`�=������%P�jb̠���O�6���s#�3�m�_B��Ϛ�F��x��'{ �����]��3���k��"��A7Z	&�d<#�^�<�S�y�(���$4�6�����[n��.bX�qA8nI� g�ɓ>7�+��Ζ�HQI�<�}3Yإ�29�r߸�+��#��LDv~��l#�n�a��a�}�h�k9���� �R{����ڋ�qP7�-����(Gc� �lTC<@�7<$��v����\�L���߲B��|_��]h�\��n9/�w���Yʮ��>���������4re;�T�V��6�2�5=kb �I����l�E=!ܳA�>G���c�AE��Aک����6�2��
T��c�<�}�=A�;��YxP�o�!����/���=C�6��{
���?�;SC'�C��r�0�*f>�K� �������R�2r�!<��MK߬2 ��nA/v�Z�N��q��k�����^̴ṷ�k�#Cs�2���ʁ��`����}\�GuX�S2$�����+�z���&�?�6�+	�KN��'�#�����?�w�!���o3`���n2C�𘿳�p=B4�p �1K��T�&��ƫ-�޼&��x�BX-ͽQ����φ�yo��`�$Wd"�k=ڵ9�m�o쓩�Y�9L�6��/�.���=Á�A���0Տ�L�|!B��&qS���r��ݤ��w	�����b|q��@{z������V�$A����ҫ�����]���tn��1V�#���~ʁ��8�g4��/��������g�f{l("�25D����k��N�y����~���ܕ�$�m��^ί70ZN�s��8y�lD�����!;��7��/ڐ�2�(��!o�H�S��H÷;�}�S�#��|����k �Υ3��Y��dn'zBCkc;5�ۖ�APܼ�A%%�q2M�z�A�һb�z������-7���FD��sB��g�j�����>߃P��Fʠg�D���O�@fiK��3��n�����{��.�	z�E��0�#{�A�L2.=%�n���(�9��s�.C��D���ӭ���)�j���x�NW=�A2~��
��v�9���ŷb�`x��O�`��.��h�Q.<�.�W�pю�������ǒQ �]՚���
�C*�����C����>L�d�W�[p��I띣bR������ ]�|�E�5�R
�0ㄽ��&�� ��.z4f��H!$�L�J>�����k�?^�(�%�ܴB��FJ�����|lD��Qf"[/����+����*��>B����?2��@�(�Zp[G�/��&$��R�U�����Kq8f��B����'��|+�֛�m$Tm�޴�N|M/����SI|����K�|�x4�6ړJ��M��C�N��g�i�2�5�34�i��� �������K�,L���? P&�]nmI\��#[����ut������W.�zķ�׈˞��F�z3\[�%���Y�����^˯��qDGP#��Y� �����C�H�4�{7�+p��y
~a:�$bW�u�O�+�)Y-M�s �WYwʜ{�;?	gNp#��ܥtN;;���[	�V\�O��jv��^�gӏ�4,��lE˨b�DM����YU�V	2���5J�n��Һ�S8j%d�w!%�ւ�PgV�0w��bWk���J �n��Kgc|���ڲ��Ĕ����Iѝ,砭�醭*�e���%0'P|ە�ׁ�y�H��7���c�:0sz�3q)�]�_%#_��o(kDm֩v�u����̮�:L�m�7_��N;���&��EA<�p?FnQ0���_��zá1�}M��\��<^�pv/�H���l��x-�济X�k|����$��Qt�m�Z�W��O�_��+w�)�dR]���6Z��W�sW��e��"Y���H��)��y�S��ԋ� ��+�A��_b_Zp��D]T+Q�N��}n��@�?��J�Y��P�߽G���f�;���D��0R����7o'�p��ϋB�8��1�ּ�mLe����
��u��8�p��v��g��P+����5e�S�j[��O�|x0�j/m�-F%�I�	KN�3X�4�;���c��1:�yv��;�e�? �H��xH�ɐ�����_�[ӛ��G)c��G��-Uo��nn�����{&��<���@�4O4-��AN��R�i&� ߥ�l�X�����#.��_�$&��=;Aܢ?FUh�5v��ʾ��*<e�l��3!��8�������"?����@�f����(�gq$]O���"d&g�u��Kdp�Hj�'ܰލun�?�r2��b8���j��y���2�CXus���yL�ɔ�N�K2+�>Acʙ�X�E��d����j�Hʑ�Y�^NaDUJռ�`[��x������}�q�Ŋ@���$�Ʃ�T"׈��q5𴘱U?D�ډ5�X{���]�G2����yT�z�xޠt,��ϰ]d����au��+�0�g�`xQ�e�#���e�`��M���Z:��z��k-[���vI�4����b�J�(ˉ�����"���1./5s��+J�Z!y��2�5hS.�@�,g� _�޴55u�s�U��^"@�d�f�S`՟�?��Gֳ��\����Ɔ���T ��������(}��N�Pu�g�"|������VP۵EM�k���@@�@����?�����]8�Si�ZS�]0��yz͍3�J-���[�O<� ���.�j�
�o���C�o��~_��B$�۫�����L�XЫ]���j.�!W(��-p��|�@�|��%"X��엤t���e���%?ع4�7�fN��As���4�v C��AA}r�L2�lM�ǰW?����0���`�Ω�e�)�S�JYL�Ky�ds�c_�)[���E
㹱�G�<���3�������ybgP
(��{��s������酺@�#��G�S]�ϔ�jX�o�e�o�H�x߫�����]�Kj6j��,�K�O)yW��-�� ��[�F{�&�ؕ����	�,C.r�ˌs�_�	b�!d�&��X��5��i�n��z�ԙŵt�����Ҝ.�D$ۍ���2R��Y��kM���5��(�p��+�-��.�.���������w|NȰ.�xT�����y�AڝP��ෘ����rT�9�U�hE>�8^1SfK�M�Q�A�
G
�9"��Qe�������D�FU�	[������$��uwG3#��>�#��Y��H�O�w�y��8SD=283��y2�r]u^�c"5~���#9e#S�5dI�گ���P7D�o�'?=�y�2T�8�n��sJ�{�$JKT�<Se}�U3��i��oe��࿞}�{\�5�a��0:L8�9S��6n�������p���p��a@O�7m��~���X���U�^��E���0d�tL�d~�U�������ʓ���1֝*�����du�F�J��!I��<u�Y������G������͢βB���r��m06C9o"�nƟyz�#��bi�,�J�s�8��D��Uã,�l��<Y��ց�f��@�3�u�w��+0ZJ4*@�R�9v���ϧ�Q�gz�_��U�;��z�����#��/U}*-��l1}�#��t"�ߦ�I��~�U��[�Qt3����Y*��9�(~��1{�.\���>��CR�1��ũ��`�9�**�,zk�w�A��c��_���@Q�ښ��g�[n�g1)̀�f�OS8�ރ�F�b�$��(�E��51�ζ%��1K��q�<w�r��6���J��?b�4��;�N҈Ux ��|�U��|lh�J6@Ca?SK��O�?^�c�-f2ҶπǖFO_aQ��[ �_�����y ��g5���<�;��B�$�pL*�	 F�H��F{H�f�q��D�mw��kx�]�I�My[p��K�d���mV5m��p+���`���N�ğ�-6���}p��{���� �����CVs�׵L���Ak�!$ӫ��<k+J���5�&Ad�C�8Ȝ������}B�8�p�pv�}���Y�0���۽fDD 
f��ѣ*%�����C�y��.p¬�N�m�B+��L��f��ΫJ��_�@��~\܅XMVw�V�nAx�g�"���<*�����Άh�갧r��EԬ�*�������Z��k�ȹݮi��aȌ�*qs}���oc_��OC�`z�G��ˍ���	�`ؽɶ�5��n~U��Ӯ��HVg�������r���͍RF����nhT�x*��CB-�G]��}���'����2��d-�?�Ĺ��G0_��qB�~|sH�U>{zk��!�i�e��7��SpAD-����Id��9�A�'�����]EѸ�+i�����2A<��ſ~c6��nMzD�''��בe,iL��O�Ac�5������4� m ��%��:��OC	2�Y) ��XiJ��kh�7w�i�"�'&��N:��؛��:��y�� < �X,G�L���@࡯E/A��Gh�_���� �������v`��)��1tr�����"� �K�,��m�� ��͉�岃}�DISLxQ@E�dH��75��+���g5n_�����b��;^�������)�y9]�f3�o�Ş��7
Dg���@��ϻ�Sϕ?@����D@�[n
Mg B���v��2 ����5��Q��q,�24Q�;.=�s�����g3V�,~�ݠ-�����,b�������n5�R-u7���F��cE�I>F_�κ}$�$�ˏ}��2���M=�3�)8�E<_�E��9��؎@`#«�||+��(��i��6#�����d¶h����B�7�,�������(�X�*۸z�ra�����	f���f�L2�ڰ����}��V�ėXi�Psj�s���Gl� ��.�zN��7��@]�q�R?��'�[������x��>`UA]����g�����k�uC=C_�`5��o��R�����QP�z#�b�R$0���a�ć8�4�(�}�F:�@�q�7��/:@�0ڗM�M�F�� �O$�x�1$J�k?�	@�s��x�*Mӹ��e3,"zb!3kY}����9^����V5��o��A��7v�X�m:P��_�t�tvPM5�X~�W�g��@s�6=-�>ιX-�A����Z�%��F�f籼�������C�9��"s�1ɇ;��x���BZ�o-Tr��s����H���_�E����Tz<�&�D]��%��l"�4���p*��ou�K�Y�#WU&�����m����$ �����"=��cٳ~�|�-(�vٲp�"6�'���|����-�
���=��}��Eߩ����v��be�`uZ��B��r�'8؀�!Q�F���+a�g�Ņ:Rd�j������c��T���St^��I��O�����Oؽ'8���x����F�E�t��fh�����:�#Љ�4�sv,��������gj�rS?�K�'n�	֭Y��9Rb�x������>��'0z�uui�G<e@/��:$r����g�	�d��VV��Z#���%c=k۾ި�����Gڵ��ȘJ�H�{A���:.�1�8���x��93k��j]�9�~[��~z��cu��O�p�'8[w�����Ѹ���M����\	��D�CQr�[��4�|Q�!.��@^�]P�'���b���9:�(x���'Dv�{����Zq�6YU��y�׽	�C\�/�ly���T:P.��BF)��^��tjA�х�a�r���'X��I�'S��<���'U#�gbX�eF�䞜q������տ;T��[Y�Ozr�h~�=p�I���#�ܠ�~l���#��Q1�&��R� ����ۭ﹎U��˱"ٜG(�}S�P̒�,������P<3���i�&��-4����)D����lm�.��W=�!�uZJ���M8��۰;��O�Q��W�ԷMaُl�0�����y��E��g��4�4\��~�ŧj^E=N�d[)UsN5���-k��ݥ�q6�����M�T�QF���C19*#e����{<��bUQ@��]��(q��!�(Wf��Ϲ���p`#���l�1�n^�Z?��HܙlKvr�9�wz*}�o�c� Z�蹽3X4[TQ���.�Ru�C�#.�b����+Lx �y>�A����=�=���7x��)��E�~���(=@Ԗ��@�X��A �ul�4�l7����4N?�w�On�Vz�ݘ���I��Yyi�!���ib6��Z�jJ/Ǝ�c�_�"�B�m���~��p8�C?V��q��?�mfϝ�f#¬�B=��`:��J�\�lLl�-m_�pg�V��ʶ���ȉ����#B��gg���?)�>��S�kO��<�5h����S �*�C�į:Pg�"������t�s���������vuDO��z=�"�P*�;]�"�5��� Yhb�.���)N���a ��ld�R���7�T�Re��]��g�Xe�D@���I�@�a�����@���5�;KU��6�6�Gd�$����h��ޝ�3h{Νh�6j%a���	������T�cF�k����
��4�i.l�ٮ�"~HN`����/>�%C+l�����!B����$�t�5h;�y�/G0�V���IiI��������� �� *�I)+el�q.�� U��N�V�f��/v� Y�X�&@]�J+!o�tV�p�b�<��9�Ȱ`-�*�"ݿ�y�9�O�}$��ׂҨ��o�HY����џx�Q�1%���~pi��U�3e^Hp�i�����LmB�aa�Jd�9v;9��`���Q�@�4ŧ������Ι�ߕ\�5�{(R��ގ�D�,3�d���Xj�+����i�'�uGr����DH��9�U��3�bi��.^���s��¿<�\�"�׷˟ZI�P(�c���Ee��>��u�T�p��;��z�U�d��� ���7����������L�4s�mJ�<�(&\L�pS�9k� 1`��/tLu�ؤ��+>�)�m?�	�j��,Wm�/`���3aU�����T�}d��(%_��f�w&wۛO�	 ��T�d�)a��� �A�Ԉc���1���, ��,㹅\\���o[���v��]M<�����*�7n��.g�i���u�G�d�����vN�?q�`��{�l
Ɲh+�ȏ�c�F����=�D5&ֺ9�cF�ȫ������"�%[I��}���7&�:�j�_s����pt?h��K{LmZox��̨G-<n.	ZS�6�Y��I�y�TL��Q�r�h[�"�k ��-��Ha>t�D1��g�Y?tXʸ��S��-{�
ա���ǡ���Gs��*@n���O�+��z�1�X�{p���O������e�kL
��Iy���G���I�4=Qy~Z9r^{L�e?[�\�Bkz���,߯��/�X�W��p��0#%ҁ%�/1�˄�	8^��W�p-5���}(�`[y��]I�4RDy`�J/��,�N��-yG�.���Kn��v\��aR��$F\9����cZq��)������E9��<hH�ap:#�� �B�2k��%�6���:�Yh�
�J�{H4�9|�w�kfL�����aކ���ޒ�,W�	����M'崀2x+,8f����@�C�/�h�}d�(���[�9�~G��'�b�*]�R��o!b�\��=�O��l�J6J���-����h|�)3D"�II��V<�܉z��\C��ڧGBY嶮�A7:��	�V�wJu�͝����D���R<5-'�t�{��z�v�]Q �j���Nh��?�hi��ѓF�[jL*��5#�W��f}
��Z���� ����(�#�P l�� -O���(��<��}ч���ߒ���ψT�Z�ˏylNa0��$"�N�뷳�b��:��q��	N�-Yq�\}ۮ7,t�糣V�J�S�������Ǹ�$A&��4����������YL[�(����v������/�d�GjI�����%�z�%��&�A:}��rp�H;�7�+љ�)�OS�-Ů4�>S������+K�u�C�{�}@؋��i�aQ��]/'��tÜ3Y�2$?���J%cp�U06 ⅎ<��=+�yN]p�w�"0@-���:;g����&�/ӌ0��=�/{/ۄM�J�ŕT���e�Vn]·�%�h�����hV��p��\[�>.= �g�|Y&�N>�rr[��j`����}������g�+]�s��;���ų4���R�%�m�E���S%�N��:��a�h5�rʜt˛�q�Ȩ�-d̛%�z��YFcT�d���!|3�$CB��Ȟ�)	xnkƌ�����->��v����4��v2��=�����cy���Ob�fC�#<8_U�o?��� �0�p>%�'�����܂�^*�0`'�g�PI��(M�"����
9��h�����gX�B�V��H�Xz ��eQ	Ύ���nK�TZ�a��&Zo���Z=j��:x�~|�����H�8�bV�TH9�s*�L�NLd]B�x���n������$�k��-�}$�g�yh*?������0�����Н���w�4��o$?2�J�*��	+D��r�����F��sM,���K-�k�0K��L+�d}�uGz�����8EK^K�����1V���Wa���<[Vh��qJ�l��"Ɋ�-M����\���m^~��h�ü���{�'8�g������y��(�;��7������I��OP2�i�x=��EA6�?�x�	j@X�h�j\���JV�f�J	�N�J���g}�H��^f �x'z��5h`e@��_��)b��οi���!��E脢*������@7��9y<��ԾW;���$�-z��͉�ς��b�F���TI�EL����tW�?��ѿ�	��/��,�Gȫݗ���ٖ���������-�X�2]_?AG�� ���S�w4�������������-D�}٣�Ӻp
�j�E�ODgg�6(ӄ�9۲bd���|��9�ul�%"]�ۏ�� �UY&��F��f�w�ߟ&jo
���n��5o?A�Y'��
��:��ÔVf�&vqEK�K4���^��4_�����.^�X�����*������C�_;m���hs���\3V�f�p��Ag��'���ݪy������?�樫����E̓9���&��
�_e�PagRRВjW�'���WЗ�j�a ��U�x���� S�7N�rm��!!>���ie����O����3$݃48)���g>)扡b�SkfA��E1����ɝ��*f2=^|�2U��p����?�Z6�g�Q��*r�T�6�I�]�?�@�W��1�
�W�}>o�@J�_�.��3��8u?}�Ʊ�8VbҌrN�k<*�-v�@��[��X{9����D4ttu��dF��f�@�_��Z$M�ړ�9݃u0�x����w��*m�����k���r��`�%?���է[gU�x��)+�ٙ�g��`7f�Ap���@��l��J| ���ʝi��m�0y��j��v���-�����U��;�R,��4�j̡�z.?�}��+�TMk)����Ge�`�v�v�2x������8Z��&T��W��`����NgBi`�D6D���
��E�;8קCjE ����Ө�br�!U!��#�{�Zƻ
���u�h����q���ǫ��<�������Ff���\]Vz̹�d��6�>�N� �V�(`��U���b�9"tu"ǣ���[x �c��U+����k*}{��(�'޼VC�[āG��=�;"$�n_\���@ױ�ޓ�K���Ek(q���!����썞����g��,�5�0�@tN���9X߄[XS�02�f؅\�W����͂H�٩�M��:a��Y!=�ߙ��?Pd ݰ��3�u�{=Ut��	���1�˿�i�憼;�<F�aN}�FS�K�C���	�m�װLi4��A��o����ʗhES0���c+��n�uH�\`�����N7�<�p���z�0�&k��.}~W��&�[�ۆ3��p�sH�$�_Vu�O' �5��h��lR!p�m�e����6I�QYg�3P�J�����}�B�1��D���kʳ�8ˉ�P��^�
�Q%,� ?��~�Ӥ��`&XY �f0���d��%V��:�-�ɿgFRK�#1���M��q:0������5�O����0���޺4Z	���z��)!�0.�Z^�cn��m�Xr�v�2��Y���JvLi#&�6�.��$z������n��e�w�^�XF�c�W�x������ �����^���g��`��R��X�e����P��J]�Ȅӿ�`f��i�m�TMI!�Fĕߔ�Զ�հ:���t:/3	�f�8��+,a�OL�'�/9��h��I���C��ʝ(h-���h:��.�FP���wTr��/�*5!�q����C&3��r��D����%���i
&�cn��G�y��Zg����#´�ڙ��?�V��h3!cat��8�.͏����`�e�3@���{�1��D7{����������<á�	�v�"܊�W�(�L���Mbn���Vx�*�S3�O�t�~_E�~�X`tU}�w+W̷�Dr�5����Z�~Y��D�y�����R�q$�MH�Ó�$�Cɮ���%'i�ܝ�⑝��e�Z�v <���x�0��aBW���c�=	�����j�9�`�i�A��q�Vh����e�6����	�����Cgxu1HF���Z�"��<�quf�c�h�F��1��"�-X��S����1{��=c�"�\�mїl�x���$��Y7Y��`�q~B��B�NѤ/C��ؼ�h'1��6"ƽ�|��3�� �s�¨�@(Ճ�I96�,�T��옋g��q���A����6�����Y\�z��)�⯥GnG�n�eR��qd�W�jm����K"��f�tB'���TXwt��R<1�T��4'�N��gE�]�&q{b��|%�%9�%\l�o��x���a7d��Z֏�"�3k�kl����(Bףy9��}
��������I�.������>�i@۹�N���Kj�p����N��gFy�Ѥ�YT����1��M3/(:e:�I~�e�s登���5�8�/c� �LJ�/��j��a�d�8.�f�����G�����UX_��,i'g��k�tRgb󘧏������Q��f6�.!+�{���ϧ0�_���l�H�ٌ�&:�W�K<��c�e�'l }�s�l�譅�-�^�n@�
�`�2����2�3��z&��Z�L�w�]j(��V�='2�"�=M����Zp�ڼi�/��iݬ�����QϞ�{���:�6zVKc*��i�չ~�����Z�B��3���I\��G�К� �?_������H�`�7��G��=3f��K��J8-*r�
������}y`,�͑�'��ǋ0S9;X���n�c8�Bz�b܆m~ny|$�>�xs��?ܻز��Ɏ�>����ښY1���.~%i�@�UK/v����ds�(AP>�H2\O���om�3n��H�`e�Eh��/K��W*�71�Ŗ�2��#q&PQ�B�Xf��eI~<5���_y�5���`]hvҞ#߭?�iٚ6G(J�`v��m��d���{���(Ca��_���V�����~7Ʃ�ǈ6��� ��S�)�;H�P�$�iGp��C��w#�A
&�E�/6��'�7lS�-���Lv>\�t����_�����k�UJ����~��D��:۶�`q1a���0R'"
'��@ ����
��mR�NfFqh'?���8�S�1yJU})� �ְ!f�nM�h�s�=� �X�m�V:����c���⿶eg�>�}W/�v/�B{�z�,Ԡ*�Y��{�*��� _ �q��\,|A�wmL�p�]�K,.�鹛�#�S�-I�營"r`~g���F;t�Ss; feoTWc��2k>��b���lPDF�1W�������j��S��ky#�ҫ�*{��
���/��2�Gm�v���	�rg�A[�rsus����To��^�v�2�I���!?B��+%��])W�ا�OD_p����n��:_++f�����ϸ�m�Iѓi�,��I���Fk�I��~)�����.�]�z*���d�p3�K¡gb�^X{���x��ze�f�񻲔�"�Tt��d3c�Mh"x����aڊ!�RZ�<B�-b����d�5�ܤ�Ⱦ���b��vut)�=�A�[G�z�F�Wwv��_w"-A{|��)��Q[g<��{k�͗�@{c�=�1�*6�*ń�� u�F&�b�&���R��1Ĥ���aa��؟�73����KȁM��0~��*���W��O�-#i����4&�[l�q`PԴ �m�����v��:����8���g�u��s�G�Zd2��.��r�JP���MMS"��"%)�;`8\2Rw�<�,<TX�R}k� 7P
�{Rq�o}H:�?��(>��|��Χ*?���?��H�(n�ר�F�'���^ɪt�����s���{�+�k����:B$���Y�lh���#V���D����u�֨��qR\!��w�"�W#PM��t�L(�ȏ��|��W�ޖ��>{��Dǅ{���:"1���RƇ@":@W���[�5�&*��r�qv&�+�����3.^}�����;��-�����8��� M����}vd�Qy�U�٠�ŗZDB��&r^�d#vz��P�}mF~QK���Z���D�������6���]R�Ȁ/���6����A��L�Dr3O^}S���nZa^G6<j�����r��3�%�����ɻ��T!�`�q8�9�[�/x���L�WP5,��k����A�N�o$�|�*g��9z�Z���ܕd5n� ϥ�Y���.��k��l����M�)�y,��+y����6Rj;Q���%����C�j�������S�c@aDgO/Q���1p��5�o�S �y .�@��f՝O�C��������������	0x>��?�����䬚;Nظ�^�R��o�,�kѕ��
�ֆ$�[��Q�h@hl܉�Y&�U�έ������������%�g%0~�v�/8�/(2.v��g�C~�N,�,bղ���({f�I��Y�~��(�7VYU
;�&���#_���E���0S�>���i9�҉@F��P&�#rqo���ivl�hSoK0εx�g�g>\1Zs-���E7��X\j��S�N�Nn��̌ld��^��L9�ǻ��v���!�PN��͙�Vwd�5N���fy*��s�,$6�ؕ��wlKt^�������vi�-�-�2�%{a{������9|��AH�aX�o�A��JR�N������ ��vϽ�@�XM��W�.S�,��2w=�$�N�r-D[�Њ�Bq�4e��ǝ}.�cL�V墂�R�F��-ġ�μ�����	��n���������)�8ls^۞R�z�9`�������vH���s�[��t����>*��}��ok�!�>���Jp�8u���%�6����#'��0�tb:0�v�ZLWt� �m$�M��Y�؃�^��a#e�Y%���iX����Z�gE�������m0�᥸!�<
����0e�D��}S��qjag	ŉ����?�BV�4V���2ǵ�ҹ����{�4Eg�Mp��]���.ҟ�"ts���\G���L&��_� �߫b�[{��&�5���@�g�+w#'��z?���O��ͅy��+������"�ot�����;@M��L���:"A���(���ޘN!�M�V�����M�s�L��΁�G6��H�.��s�H>2?�Wn;pd��pR^����D��3HCyt��d;�CXQQ�־����/O� גZ����ʃ,�L&�;D��DhZ���G�s+!����ȼIA�$�m6���b�Ȁ�p��w�RAHß'�Р�u��#�S�̍�"�L�1xH`DQ}��l,�ՠb�5��*v>���
���cb�F��T�r/r��7��Q����&sF0}�����hlH��E?�h�cد{�����}�J	���Қ5$ই������`y�� �V�f2�6v�q')9VѥL��GcJo����r����Y��p�fz�
�ӡ���*���R�rZo�hC]~΅k���wF+wf�rB����hs�F�>θ��@#}M�p��2��>�P	�	��R������~gC{tD�s��5C�b'P���I�͘�������%�WI�������|��`��7ݻ��k�6逪<I�.��/�2�a1��[)0)�E��E��DeK·��y�	xE|��č���F8d*��:H��at,9,/^R8#��4�q0�%űf��:����?�4&��9�_�y��1ׇ
"�b�nq<�	�Γ8��}[p��O�m��.�5*��h�&�����|���wVP����%��
3���3������
�T�p,���K��gG��8����@v� @�5�O�{ܾ�Ξ<��⫩v��Y������A~)c��&/UЏ�w��[��1\䠙�=b-��@��y�7�׋?�e�*͎7��PT��#5�v#z��W�Mh�y�8k�0��V'_;�_\~s�p4-���)Sg�0�W����cL��d��fbmm�f�mA���.@����$��.�nir��+'d����������|P8�R����;���栅A����eF�
��o3����eӲ��L��C�m�pa���x�:6�"r�6�SC�:K���́���x��_	��}(�C��X.�u���c��ޢD���o�ţ���>������iq�SA�ل�v�԰^��z�Q���ð��R&2ldʨ>���;gR�k��?-��F̣O�h�i���]&�l��.W�xQ���n\/<�8���7��N�J��X�wY����'̱�(�e��ܞC0c�V}(9�M��D+��El����a�ͯ?X�����
��|p��	]��ʉ����w�x��@�Tw@W��2y/S��C�*3�N�-��h�uY�P��miު� �@�V���gA���O�x#������o���Q�BR���	Q��Og�穯��;�J�Ꞷ�B����o�*���C'�D�� �)��/ǲW�*_`���<ղ>�x��-�Y���~݂��T,�����t��@�4[ȟ zw�hk㫀���J��p���Z\#�bX��4E�q�d@9�!#j��_q@&�ZŌ�۵̀��F�9�*�&W��ر2�ۘ������&��5O	n��=���SΌ�)�6zc�kP�����㴈,$�	��P%�線a�i�{L�����:j���.x楤4��<���W�a&��Iښ�1�X�`Бz*�i��w9�Q�f@�%�ޮ�z^܎�M|?���/����̅�����X�|~�&�. ���6@��������U�،�[Mf_�p�Zm�P;��9�K)M\���!�td,�Pn�s�<�g�<I`w`z��5�*N	��I�8��T�hJ�U�H�V�~�"D��%�~��{-�� �Q;2��/�脡�S:�Ɨx-3��;�������&��&�s����Q���v.��.�Z����%x+T�@�tL�q�W��iqB��pZ�(�<~�s�`���+�Tw���������ͥ�SBr�gwe� �[��x1A�T帪F��M�B��<7��)7Õc8n�\n���!u!���ܞ��Թh�� (��v~��r��Drp�/�.J%����H.;���&�%��\��Y3�$�A���]�5�t0�F!$�׊uf*����r�2 ��H���qs�������?�{4���F��f�5m�!���3ll��&���g!���;qi{U�nz>,��b��Nj�/<�� y�o��0�7��ˆY�\?[����"Z��[^�%%�=[퍧l�G���A�����k����,��ˑX���Q!fM��M ;|��DG��M�~��w�Djj�^��IK^�O}���S��F�2C�|��#�_�B%w�V��7˖��yZ_�A>B���p�WE�wz���"4h��>Ɠ������v��1�̈́i�E�&�I��r����rN���]�U$6[6݉�Ȳ/­��h]��$o��������E^ㄒ���Z'�ʸ��c��������m���ڟau�|7qt0��%3c������Ȳ<B��J��BbD_Lj�Iz���;/꜆TPL�U�'�k���|Qī�r;!�5�{��4o6������Nb��,g���3��O��γ��"��Z�]`%���[["����q���J����d���5Nӂ2s�O�Ͽ�<�J2��5g6:�?�ڜ�$�x��c�%Z%��ݯ����}ee;q����Y�l�E�5���ϮK��0i���T��x�4����aQ��@k0�4
��*h�s: ?C���1G���Ic����]��(����A�����䇟���jf~Q��$N�G�mH��@�xH*�����ը{�`���R�]�R��8���B��
�� �:�����M��k���h�@^ם13�06��|�rH�з072J�_υ�k�j$�/'��e����'	�y�\dLr*�A���y����p��D_@66�;��W
����%gR�ԒB!�4����H����"ph�:X	�Th&mf[��q��f({'T#��#��yt��
��W�LiP-���T�s8��0�����^�ۺ�V��#K�ei�\�\�������e	��
�>�Y�,J���7���Z*nc�0v_��!Là��%=R�N��5qوG�!�]���]���9Ğ���+G�?B\3� �	�����{k4{/ʥ�`+�f�����Ga|z�ÿ/�X`�(5�l>:���f"��;I�����6��s|_o���^��HvL��Q�G\�	�G-c��m��H�6�J����t��=�/e���`�XD7�T4��%+�B � c/Wf��o=o�C��	�[X�u[���9$��V�׼bv�0�M��KZO|P����g��ܲ���B�Q��s�4��or�
�+����EZ�h����:aGo7�A����݁@�`�[5@\0"%��{Bܓ̕�^�4Or-9/�g�VJ�AA�a��yO�n�~QCzx,#�0��F�5A	0�}��(U���m|^,�^2`[q��*�q�^�0�O����Cc2�FCs�Z���JO>!l�۠�A��3~q����x&D��pi�S�q\)����=��GT�i�M�6Uzp��?2�Pq�������+�I1o�
�}��H��+cVe�`B�s);�R=}Z iE�!�Ĥ6�l�U���)�D:�g�?X�^F��4놋��H����� �7ʔ|�=8�!�������f0y�p{i�XѴ��@�BY�)��x:X���{=��Tw�F���/�f)���/� f=�w���6��ڒlS���m��p�����Ѥb��_@��:(Mf�q�u ��lWC�\hEb����u����-�����!���r����^�rg
��?��9o�0�](�Kf�j����3)N%CR" .���T�&��N��O�����J��W���(Ĵ���@f �g��y�Br����Y-2zM�u��Yb�Ӣ=s��k��L���n�"�j�%Esi�y�D ����ſ�[�*��YN�����K��<(�֞[��jUϤ"%8&ϫ��kB��{P~���������"^���8N����9��kOtq�ێ��Ƅ�2�9�p���]�����iv ��E��OjŽ�Lu����G��\Έ%!T��j�:
�杺����3|�D0*���4���)�=�b�{+�u*�	Ȱ�˫Q����N��FOV��џ�6�fh��9�+Ju8*>���<"��d>�_ �*��x >�0��F6��MYh��*����uU���� 7��r�#�d�2KOu�3[@����4��4���R��i;0���}	�>${Ե��)���ꬑ]9�Zk�������ؚf����: $]�gb�x��rȏrs9}ޝ�*������7� V�������k�S��z>�R:�3�S/b��Ԕm�DI'G�mt�e۽J�B��6��~�+��ah��
�i탸�Y��*���!�[O#a+��#�~��˻���c� ��t�+����B�G���w	�+�0��B��7,�ݍ��8��r��#v�!s��sPC��ccG#.���n`(����d@���O��`��|P]ۉF�:ti�a�$��9tM����_#%�~=5�iW��lWU��g�ˎk7)����6WҬ$����	�����>����bQb���yl��%�2����M�%8-9���qu
�>�L^~`��i���𺞵Yt=��=J��h��e_3�Q����"�~LR��R}����Z��)B&�5�Y}絝9[d��V<ͧO%|��L�xz��G����p$�I�m��uf�3~��_��м^:�ǽ,���C�����i�|�҅�]��`����_�i�znсork���P6��é hp�h�{��eb#fֵ�j'�lՉ�fwL�g���c����\�y&�����_Ps�����y��ll?jK�Z	�;I���,o��4���!  K�}kk�6���Շ]n��v{ �Yy�v��-〧3n�B͜1��Ry���,�	�V�-� �Hs\ZI�na�Zy�n�ԇwQ�."KA�d�����H�׾Y~����%Ox�A�UН��E,͙���t����c��U��}bس����9�O�L[i�g�X�.��aր����!Be�`ӭKoq���$���Ts[nr�n��⧻�n�Ȍ�AT$�܉�4L��¿��^7^��D��A���u*����K%1�5���o#j���oL?�����:���m��m����g�t���'1��(���ͧXN͉j�����%�c�8�ǲi������M���lP#��	R��)����tQ3a^,٠�|}gg��r�D��{�q����&�ע�Zl�I%G�?�?52J����r��6&��O��P��,]��x��ɯt��{`���$��d!�Z�,ܢ��a<.%A�x��of�����݋40�5(硱�:<|� e[���xY�bL� ��42*�_	����i�H[Wd]^��c@��$HY��NЏ2b�)�m�W�#1X��a����u a5n˹IؕY.����{y{�;�4�:ԛ��y��JF�D��qj].� Z��-n+�rD Q�^Hk�~W���R��������{�t�q*�m�&��ܚ:"�6�k�����xEO4�]1l6�X1H\$Aw�Մ0��r�����=���/e}nm��u��M�E<J�s{��k�/-�K��G+�s�	x���*q�D�i_�K�嫹�f;=	2V[��:ZE�Mv��xh�������ߊ>F���#� �GOҢ�f�ֹ�@�. �+��e;�z�?h'�c���Wzh�7��Ja�����B6[1O��I��lɗ�������B>V�z��r���c�V8��L+=�'y��?�aG/$ƝAx�w�{:�Iw>R����������X!�$5��'�	gvy��P8빐P��cC����K��pU�p���%��oXC�M�iΧdy�9p�E�|T�<ɝj���|b� '��$�1ˎVr ����qqm�Ip7g;Kb&f���Cz���\���F-�&.q8^\�W��;"6;F:$�Vc�]���k�s/�څc*�ڲ��h0G��_��*Ej[���T����.r�'v��J}r>��\���d����iu7튜��W&�
e��G���QĤe�;Տ��/o�<b�U���	=�&�1Su�Ĳ�p�t�0��m]Q�M��o�q�MOk����F4(�����O�E���T'�b4j��	~���?5��;�8!��H��g����x�S��ӹ���#��O��YX�@���	�l��`[���:q��x�q��8@���]�{�-Y�Q��K�+���8�q�OKF�f�A��������d�^0����1��7 ��g��f�$���N˗n]�wr���ɌP�/�-��,s0�p��ǘ�MB���v;���/|5��V}�ڳ��a|SM=_��ϐ�|f&I��I�EF�7H2�p�YּP����d���uB��"�6v&���H'OP�$��Z��τKRd��q_O��yR�������>k��N��U!j�r�yf��"��a?���P:n.�"ن�=<w�Q�7���<�M.��� �5X�͗����u����1ka�Z�K��|�����*��E����ͭ�W��%�� �C�A�*��X�2�}^2���f�laa���3���Ϩ.��#1�;���:;����g�#��W�B��mvJ�&��ѧ$]51�&B�|�ؙ�r~�u �T��^�ƿo��7�\|Ҟ�Re�֍�~*q�{��8�h|�_��Oe�(����NS�po�)5�}��~A37��2G~�<�W��wd�����i�3�q�u��$�(��]�-W"*.V
�%�k��%n/�jx�'r9f{x0�D襇fH��{���,����
����h���r���%�B�37ǆ�VJ�W�F���O>�2׎ԥ�<H��᎝�45N�.Hc�&i��?���*�Dcl�=0��3�_Yc�٨�g=�;�h�$Ӟ9~����N�~5�ހ�^q���jr�U{�3�O�2W�!L�/#�p�J;P�~Q�i6�N��9��+5#�����ek��/�%�9��ވqKv�{�Knƌ[\3e�IZ�TA������y����+S�&�x�@�'Ô��̜���2(�-^���>��}HN��^1��L3,��3�n�h݀(��c��T�����q��\bgJ/q���4�yq�#���Y|�Xșy:[��M�h)��j"O9h�z���v�4�He�R.w��B�OQ�]K���(��"�I�-�Zn�������gz!�as��_}*�q��5
}%�u��Wo@�S��� Ofм�`�=��ڌfTSѳ8��}�8�
�s�N���^���b�k~D՚ ��2���,I.���P����Gܬ�T!{���^T��l��&�Ȯ^�'J3L��֕uа6>�a��4��Ws/�~�&��\�q�+x��z:�g���,=��Bl�Lұ��4�z�����ʡ8��P�5�i�=�ˎ$(�@r(ܝ�2%����'mI�5���v%����{���w����K@u���7�%�|+L�#�E_�����.@V8�2�}���hp!ew{�m)
������'��Q��&<.�ܘp���~cꍘ��䙞|&��oW؛Jv>מ��[N��NOf^�6�:��L�{r�V���Vr;,�l�����uA��E^l�kx���y�r�p���o��5'0�L�ۍ���;ނ �X!��
�)�{P ;��ĢX̏b�Ag߃]���	�!�(42aZe�H��QH�5 ��W������ܞ	���܅�K��n�\�GJO����h���IR6�_�Mr{]r�T�U B�&��z2-(Ga��%a'j�K�� ��I���0������#2o�n�s=����4Z̉���1V�J��lF��:P ����
�n�\�67��{�``y��==R���A��IS�����T�:ף+�/l���c��?9{��U0n�m7��g�k%�	�Ԥ8#z��W���$�:����sm�8��oq���P�E�kg1.��E�<�m�kD�ҙc��w-���G�$GK���6��k�6��݁��fx����UH��~��2-������}_�gW��$�ӕ���u����CH��n��E�T���y��%�����:?��f�����uF ������V�����.]�]���ZQ�xZ@��߸�*��ț���IT5 ����+��������e�:2F��%�>�����DNj7mHO���m����|�=����#�5��1���P��`{�A2fb�O���a7�'��wXv"��Z����	�w��]�DCKP��(��*e���.|�p<X>�P 6�ٹ��m�����xPlVO:
��q7�����r}��kH���?�!�V��Y�=�]�D60eu�\�}q��u�K��cc^h���7G�thEק�5�;�K��X�,��|Ұf�A�dq}�y���x��o_�C���5���|m�QC�%�,Sk�����
����*�zw���<�U$�J[H���w#L���5;����o�BW#9�x^�5�`��G�lГ4>i�jIۦ�]~h�k���a�B�*9i���:_�S���J�*ٺX�o��]���{:��u����T
�=����#�Q/`�1g./ɢ95�i)wQ�6���`����ھr*�|+�(PJ�a���������Zc�Ч=q]�@@���]�lN�itӬ���[��+���X[B���@D�Ă��o����قbC5�F��
f�樟"�as� ���n)�jT=����.}"z=�Ϊ4`w�C���=�1�X����w��Ī���Z�*�����2����PT��EQ��
TGז{�J!v�ZzhA����s�.�',�ԔI�p���5�^���;�i�m�|���c$�bJ���z��t���{
��l���E�W�P1&�O���z���dH�e���!R�C���$�U��v�=�}������-���0B��U�E���VyM5����O���4��	7�����L��8��Sf�`�t0.�7"��L���)�ꊌ��55M��ط^]n��8��$�X�h���^�t�K��v`fA2�;��6���YlB��$PeC��B}䍧!����b�\��z��L���V�ɃtD*������z3x�-.���)�IX_�7J�<�kЕ;!���~qM�6�P/���K�ƾV�Y��OF>����o��'��q��ڍ%���W�o�����9,���cSA��M���b]Ml���ߦ٣H��-fn�%U=*��{��x�GfS~@�Yo_��dc��#�/����;�<�q�<&���SB:��{�@H���u�M�,7h��̟g��YW���\$=�O�Ԣ��'Wt�f�a�fn��;[�ƊT��q����S�*J8(�Bf8+1����S
��YwO�_n�4�a	5��6���(=�q|Z��/6Xr17]��_��Y*6a��y�W,���3עք4���چ1��?D=�6*��i��3�	Uw�ޮɶ9Ɓ1�����t%�(���@�0�L��?w����GgJSЦ�y����Ɇ��˯�!�og0�7c�p�Z~3X�.)��c���vQ5z5���jch׆�ϡ}74ET��߄�+7���y���u\�p}�P�T����9��c1z.�����H��<x%���Ԙ�-�����2��k���؉�>�C�n���=2�%wV��� ����ڊL������IF�'�@0J}# )ف抆=�ֻ[w���/D�F�V�K���őa�����l|�d4M���\6��5ȼG����K3�A~�?�L�ØEeB�9����\\��~R��ަB����ü�W�ҟL��%=78)�W�����c�N�@��jy��Y&l��.'���Uy�W�uS0�95д��a�.g�eC	�ddv�մ �7EO� � {0M��[l�����_@Nn�C��^�i�;���-����r������0$�5b^T����>��E�X�x sC���u��A�:�	"����J�d
m�]H1��]�@����q� /�U����<c!�C�~�by�����B�l��L�え<�����sW�|h"��h*�l;��9�
+r	F�b*<x�q��HEˢ��B,'��@$��M�GCB��_��r�?|5u�����3,��	��FQ^Z��);����4�+r�^�>̶z�ہ����=�\W�J_�Z\[�6�1�6a��E���c��1Y����|��6�ܠZ�Ի�媮+���C��%�>= &Ʊ:��d�2��@Q� 6�B��J�v՞��V�<&���>"��'2��0���&�/+~��G)��.�~�tg�l*۟ȑWy�j�]���F N���@�M��D�p��9J�~��D��8�{:�R���sF�k�vՑ)2MI��1*�1v�� �^)�kC��Ѣ��P6�ShOٸ�dy|Zh��z���G�.eE�$�-�y�7���q���ۺ��-�[�o�;�s�%@?4�s_��?\%/�S���K��O]�/v� ��TR���Ѓ�n�x�0�S�8pN�8~3_y>�R�W_3��Yg;�ʟ�~�5�z�CvP1ta�Z	<�^��f?�Pc�N"�[�ĂUO�9<��*�ڋ�_�;Ia$�4����x���dL��5p�8�K��V\H�:m�nχI���
��yZ4{2l.EM,���R��EH[,E�ǯ�! ��(�R� ,�i���%�8�2�"���+@:uN�u���}Ԙ7������r�.TJ�/�\�7�&W����nt??�F����e���x/�MS5ZW�.�.%@
~�������U�3�X6�\����?�3�Z��ʧӄ�Q��0J����b���q�@	Ä;�KI��roJV���V6������|����U�xA;���yk��˼��]0E] >frV����e�(�"le.�T�c8��$������y'm�)WC�Ë����jg��.u���Z�|�����f������?c�
Ϲ<8`�]k!��W0n�f�L�KZKe�4B[��n���d� �*%����BZ���D�Ci
��ik�.o+k\���n���0������p�AR�z,Nn��o���<5�d�MQ�L�8.!�T_�p���{
M��A#ڪ�b`�v����ʩW��� �~�v����s{T1�Z��.��7�'�a�x׼"�D�|bÏ?�OY~�xZ� ��K�s��S<���Bp�J�.���Ċ�TҺ-p��LJ�$"�0�v�a�V�/�&8��Ep�+#������.�O��*#쥿S��}U0zN* �8��g�F��.r���YbA72 {E�w�P	���. (Gs�t0��zI��V��<.ժ����'�U��8ˈ�D�x���y�������x1/���`3/���L�@�`���򈻋�Bhd;�7Ď���}V��%�EBY�������W2����Kse�7�z�0O�Zi���!&��6G^y?��su˵aÔ�A%�ѡ�Ij�!-���X��F)�'���e�?���9��D#t	����3	]��S|�P�5E3N��4�P>`1�y!��>��d��1|���?�QIo)6�<���0�*�N{0�_��<a��ō &LC����W4�.�?0H[ ���R2�R͇��ʾ$� �L�I��x�$�/F6�Hu�d ��op��m�����yE;vNF�e|�T�Ԕ\ ����1��l�Q���Ⱦ��B�D�e��-���s_������B/��$
�g��e�^h�M.w�H����dr�ھ�P�%"�����LFJ�{��v��,t��v��ȧK�y��[�0	d��qI
Sy�ڤs;uF������_8ǁ�<����-m�P���	�UT}^����vw��3�g�vY�v��0�I�`MW�C��VD�/�{����9�,���&�$�)|E�����{ۋo��plJ���uŜY u���� ���B�]���z�(Ĺ�o�C[����N�>2�D��.�r�/�E�UqC����O��z#\\���cq�wF���3xĠ�	\g�0�q�͗M~��[���k���jAt(�Z�Nm�¸�*n��g�	�g�,F�ʝ0��ҋ5���ɮ�.y�n<��N�������[W; Qok����������.h�]`C�h��6l��4<����aDZR��W���"��o�ʞ�f��� ���QE(eE��^��p5:��l��'��rξ�q�;_���
Ō���
!���b��G��E�}v�8�O�,� � ��-k��K��w��Z9����Jg��R�G	�a��0'π�V�	�P�p��Ry~���k�pWfʑd���g��o�Ш�^ښSk�aׄ��I��$CE��G������r<9_�[��D�#ux�1��
�ⷩG4�X��0Y��)�%�ҭ/tC��r�ꐵ�$�<k��hxfn�N�1�]&�u#a���$:)"3"AٽWݺv��[�d��.�pP�d�X�#�s�l}��-���I��Ӓ_v�Y�je�O����O�i�>z}�nž<��h�317H0[>�pߙ���� �/e���B����&xO� v�����p��R_��N���y�%�T�������/rg%�d�����et�vǯ�35\�>�% "'���^$ׅ�i}�9,�\H�}d��H�M�d�$]&%�&�Ib�Go��)���r�?㐵���n*5� ��#S�w'� 	Yi���Jht};D��!�T�d�Ҝ4.�[�P3*�9ȘH�C#����-T�2*�PU��.�Q��1�D́�
��sL�@i�՗"�ъ'ʹ�?ż�3����>!����\[��{܈뎧s�$g�7��SQ�ޅZyR�>;K]~�@�GW���o�A�إ�v��u'�d����A�o���8�dFe� a�M��|���a���a~�����}�I�n�H�i.��?啠��f��#1֕�l�ԥ�x��W,���ò�_2��F%qnN�W��7K'�J�7������ty0�_ẅC4b�CZ�[�;n{r0wlup��-v�K�S<6�j��wg��_vgգ�Ʒ6�v�.�!�YQ��"�E�&�^�b����{��<t���cT�U5�ΧA��۲������tM5)\��|1`v��bM�u�F�8�Q�)�����[���K�A]�q*R*�h?{�={L�]�r�5{e�wm��*>j�;��l
�W?����"\�r">���@�cRc�����0��i=?����Q`�TǶ_� 
w��w�T���H$s
Ğ��<�!�w��O��U�ڼYo-ǿ>���&��~O�Ca�/
�*.����,�c_�\��3�b�J+� �Dc��oo*���EF2p@t��hk�O�d�p^-����?���Tȼ�Ik���b&l�h�g��t��§�;QPĲԈ�;Ӆ�,�%�n��J(ya��2��?�c��"}5c`��#`Z�=�OY����\�,b���ns�]�|jZ��p�|+k>��v�%,o4\��vTҢ�SAI�3�����k��n]9���"E=o�b�jr���W�~vwSB��P�`�d P���ޣ�	晢Ei�aC�frp�k�'+�LtV.��N5��h��>�������`����B⬽��0LX��>L�7��po.zGy��CG/���I�Y�x�]���ВN#t��/C"mj9�<�w�#�2�)��q|/	<��k�F�^τ�/��T��lU�S2�˸�	������1�l���7�sfd�5YO~�ψ���;��<�ᠰ�o^�Mn9��u^�2;�D��ٱP�4��l%p��A�	�{�ݓ]��>���<�%�F�H,���d�N�Q���5K�T�щ�W�����G���:Mo^a��D�-�4���F\��(��ٯ�a{�U�6�9�xz�,ϨTV�d��I<���M1�����GÅ6)���OW�~�w�M@�~����׃_op�V�elv�콘ܹ��=
�<�7f�~�P�,T~4,\�O���8���c!t ���D�fz��Go`9���1�k����ڌ��c���ŧ"e���x���js�-d]A��&jbZ.�]î☗���d�]�I��:����7�O9U�ӗ��9�L�:xW�x0��df�0� '���n��r�V
��5�T�6��T���o GDDqy�ŲVQ �L��:��D#�Q�(�D���P6��
��>^"���<+�_ז��}�����{j9w�2�R��_0�m>d&$�����D�
y��=�>i6M~ Yp�k�X3ʵtn��� v���_�����6�e�Z`��7\{��A���I$B��Q,�e�m(���~`T�S��t<�|�$��2qE&BY�>_�U�	�k��>V�򔐝֒aB8��2(��u���O?� (@$-�{LLqhB@m�@��L&��ؔk|��[+�R��w���>��	Qw�˪���+�)ӝ�Ϫ��r��dM�g�"A�?տAΧ��Xb�1��,�:'�w,y��J?!} q��4��axҸ>�d,|�C����L�!�*	n��)�oAU�q��5)�UG�f� ��z����d�+D�Է�����MG�y���˟8�uL�G����sS�@��ɹ�$D�D����:b֭GP������X���.N����G2��7̝V:�[�&%���U�Swϑ�KW�N�;!����^	\����#)Q&��2��BN_u��k�u�Ǉ�4a�V��S�1;�l�u��Y�!�TM�m��� �ܖ"ߛr��Ǘ<Ӄ��e�Vۭ�X~���f�A>����3�n\��ޠo�����&�n+�w�j��e�46i7��E*}�5������.��� ��p��}
&��5LP�(-��DN���t�8�D/S�pq��j8�`9[;��B�I�G���0ȝ���k��j�EI~9z#a�s<�C�F��&A(F��D !U���\5M�r����߿9e �;��uZ�srei�� ds�O>���b�iV����m���ji>4��cH�G���[6U�4 `�m���F��Ð@$�u�t=��2�*s�j��h`�Z�
DRK�N>�-���ı�N���K"������2pԘ�� r���U�t?���󼊷,�T|��~&\I��{����R0�->�����OȌb��IK�,~WJsE�C��Q��]���5
��J�Os~�*>]�W+J��<w��p�C �?��z_�Y��9��޷φ��d�E5�%�-b��1����OZ|����nSiN�)(v�.�97y�JBÔjWܪ�9��������Q8�f��ՄE�.I�.����5�9J}<�xm����@kx� ��h�o��ǡ���}��"9�*�G������d�A>nmr�;�]������Z���U��x��Rz��!�ƽ(PB�:Ꝋ Ģ	�R�K؅q9[��)I3��>TP<p�_��Zo0+J	4k��;�R��P������N�� .��#��R��M�Y��~.B5����V�vA��]��P)!b�����ڌ��so ���;���7�\��$�Y�vOö�}�+*�E��b��{y��鬻��$f9q�.� �w�S~ܫ���u�!���_D�զ�~����NwN��f���N���@;1��B�Ro������.:{��}�/�l�rc�-�:����7���Í �0y�{�xR��̑xU�<��^��U�����Hj�����G�3�,*'�����ݢ�Vj^Ƙt��C����L�<dM�082���MN����?s�t�QZ	ѽ����!}�����ȠI�u���W��[s��_D.�����-�/����X���eZߪ�Ѫ�s ��`��B�Eã�X�Rˊ5���Ǩ.b[^A��7V�A�n�G묕V��^l����\�4����^D�`�c��!� ��r� :�l����#N7�N�<�Ls�sO��jQ���"K���7QKſ��ZMn�܏.��w��B^�^^��X?b�E��2���k���d�A8�c`C�B�8�M��?0�Y��2��,���`��Ӏ�ٶ���SM/�tc�U����=`��s?E����!.?BiI��D^a������]�e�í�c��>x����t�J��\��3�k0,jֿW�D����|J=�>�!vaEf���[o�`_D�-�X�va���!�te=��M������P �7�m�T���u�e��0�Rj��\�v�P��C^� ���za-A�"��Ur!������c�I�3�W�Q��,#�T��:��'3��Ue���V�ϰ ��!��K�@�k�ԝY�)F�6d�[�Y��e�$Dw�H���/�c�ѵӾz*���`n��st'����[ s8q��V§s:Oס�)�>�Wn\��6ܯ���9�jr&#�xuX=��BԲ2�H���C)g�M����T�k%R��8�_\�,ks��G�t�#��Cr�`��S��/Q�'� ��H3e�3�k9	h�r~�fBR�J(tE�X-�e�XV��J
'TKo�ynYi��-֯O޼�:/h��EYy�Q�bʈt��!'6��v&�9�Ia�>�ü�zh<^>x�N�} pK5��b�U�v+G9�XN�Sp[��*З4T�p� �1�AVGa���Kmh��=V��8���(C�S����� �vjC��t������L�Em['#Q]�Lʺ.l�;=�r ��n��qo�oDDq�8���ne-��=	1�i���h�ƻ�d���\BoHI��
,��KS��`�������|�ޖ�L+ʬ�F�YS�d��@H�x΍)���RhQ%�@�;n9/	m'�� b'PτI�DH�v��䶨�%��X��t��Y��chE8�v�t��n �ؤ.%j���#\\(JF�tXK%+�A!�Ay��4_�Hi&`��j��տ�O�9��B�(^����G�D�"��� F޿�y��K�SD�c����Rz�O�����1H�Y��H�J(�ڳL6'�v�%C��#"��������D=�3��~�����R&m�r�e��H�������J�aͦ[��l�1��pS4���ah��7�����XD�9�5>s9�F����I����,��i�����|�1�Q7�v����i�ͱ��BMN��|�k�d[B]E�"���{6�2,8=��~q�NېLF[��,+�*�r8�B����b-.���W�^Xt���]�����K#�6�{կ��[�b�m���q>��W	jeB���#��n�-V9R+�xų�����W��M���eQK��%d%�'�w�����]�!������w.�` ͤ����O�n��j7�����3I�Y��ky�y�/�!�/���]x�w���n���4�F.@=�_��+�{������^���#�Bmf��N]�D9�h�%�ӡ�H��nؙ1�� 8�����5e9����\@�*�0�]_i��3�[�TGZ����5O��U�AC$̟Q��xޠ�;qY��ٳ2���0JG�#JE���(��d�����+��J�#�e���j�T��@� �,E���᪆��(5DXk�g����^���JJ��k�m��L���)C��TU�JP���F� j���P5xd�������L9��5@9�v2�t��icQޖ!'^Ba�D�̈́���J�[�Y��!'F�,Cݪ	�EZ��#�W��g۝}�D��(SĨϦ�b��q$H��\8zj��\9�Z0:��TaQ�VLka�����JW���1T0 0N_��g���6yc��x����	5���mzV�m��d��ڭ;]ݭ�r��|䲴kU����^?ʱ���x�Dg�P�*=����(ժ����M9�Cw^S]�6k���2=��BQo��4~B����)�&�Q�s�C˩�z�h��t#��8�km�]FM�d��,7�V����S��C:Sh3/�RF�`]V��-ߒz_B`���Y*��]�߄���A� '�S�%��_:���9n�d߃?��
�Q"����7t(�t$n"��	��R��h=\˘�����]"��lE��'��S�l��
x�]K3!:,�>�Ϥo�����������g\�/ta�b�ۘC)�:fȴѶ�q���`Q����ݕ�
���ͨ4���p�g����;j$�oݍ���]WǬ�Ǵ�gNy�J0u��^�*�ݰH!�����┱|�v���}�oκ6�+ꖹ"�cQ�����ݍ� �_�����?�����~��]Su�>�s�jJ��SV-�Q�˗�E7��\��O*Iºz�XKuy���R0��E�4�ʹ&�D��mw��z�90:�����_��)e2,�B�Oʢ���P�p���G/���bUZRrbdHR
\+ʶ�C����!�jl�ے.n\�$ۖ͐�:�B��>a�B�;5�&|�:<\;���%ɤx:�&éET�j��vG���0�P�v6Q5Ӑ!��l^a�M�Y"��F2f��9�s̩��⭊=�h����Yh��;P���T�r�W�IV�2!���X'�	7dN�����q-]a�n��,	GO-�m��`0!�z]È6��92�u"3gG� ��d��k-�t.��AGS	W�#�7F%0v�r�C�NL�*�?|툠p=H��BFq�����YF]�pu��Z���Ze�"��Ńeȍ����1nO)���c��0���)�T�<R9���gC`�pD�ᓒdZ��� $D%)峖��e�o���AGm���S�F�1�r09�]��f|�ɶ���hw0�	��Gf�#��/e\U2{��H��P>E��SL~{�0��=����Q�p��h�}4JXtA�$KF�<����mRO��q �gQ�����%�vw4ƨ���@Sơ���|��ܹ�o�9ޔ��� #�vUjuv�7S�kQ���A�F��ގ�pk�@����m9��ԭ0����g�e���H!� �[vD>r��ME�Kf
Q����٠/�$C��<����X̎2Q��'�(�\�@1�v�7�	��v|�{Mѿ����
bf�ƫ<�XA���N�8׊3Z�M��=�GdN����lS���)"�U�y1�E9/�O5y�?e��H�+��;K��=�-�A]�Z�����ު�"�
nz#C����})~a*�
m��K2�'�MDK�Ǩ�Q����zTR�h�վ�Cqf��y[�U�>��<҂�a]&f�i����a���eWg���U�&|��^�ɛȉ5�(cjE�����z��|[DT�͡b���>l�^wpӢ�>D߇q���h����eT
��Ӳd�t�UА>�'��O]	�^�㹼���L����Z͢�Dj��H�/u����B��Ŝ����S�=�$�2d�֨�@�-kZ�./�!�C����m���u&���P�z�XL*�h�2o��69o�Yy���ٺ�P��{)���*I��iOR�����d�h��/q��0�٥�%��V� �
���2M��wI�j�[�^u�}�����<�A�1�@�*	E�z8s"쀶@R��m"�+N�Yp�q,�lؕ�Oh��*#b)̨�$NY[���sQi�~}� ��aV���΢	�mϓ�
�q��y��6�sguG�g[8-���G��wԚ��]�'ԝz"{6�~(	Tg�=.S����?����)�_Eww��<ܷu�粒����RO?s�0^+�FA�;�2U�1J�ϧOm���(��Ǉ̃f��q�����^ �D��r3�Z�v��)�X*�,�kS�~�tT3/fo1Pg��:4)�g��]«�pj�Y,Vٞt_*<��-I�^M�����,!�,'��Ђ����(g������{���V�7��1|n:~~��6LL[h�?�! �"N�̡IZ=Y�ك����&6m��=�dCW���b���*9�/��Y<ZC�ԞR2�Q���V�#�R�)�l�i���P��:�^)AR�a��:��l� �c��
�$  �9�*�oוՇ���Ǟ��Ԏj�
\S����Ϙ���ch4����f/���FbnK�ilc�Ƙ`�4�A���c_>�.�]qvq�"�g\4/@S��P�#�KKLN�Na����|1�� (������X��)���]�\rz��y{}2��4ʹ��5?�B����Ayu�7d9�s��R�{3qM�~M��7��N�u�ck���7�.�Wp��A��i�?t��^�}#ٻ����b9Cv��1�d�v�*�񶄯n�ˢ��s5����2��̺�5�:ö,F�A���r]�8$sR�.~/��%#��D�e��XYHa��gm'�͙oiT���f��P��Y/$0LY�G�>�ՙ����r��J��)�.��/ZZkibҍ�m~�q��*����цD��a!�T���qK����k<�n�2(��m5�\��``��߷�T��L��x���̤��'_x�֞SЛu�M_�v;*�C[��^G��۝���/��=��i`�ɨ���葲��Ɩ��H�0iQ1��&��_���&�u��_0S\γ����G^ab㱗����p�1|ge�(<B�0�y�DYI�@���"iN��R���9R4��|��.��I/���ބ�4���(�Ih����=��� 3��3��A'�lxU'����&��c�klE(	Gi��
4��̳:�:��g���R�A�G�����
�"����g7�=�q&�`�4' �0w��lWa�U��^���	���5��ϴ�s�����AٶrU�(�y8���u
������pc����4	���ۿ/��б�i�ek�����%$h�{))���J��NA�苇88h�{�=�s��+ͩ�v�^�WߐmZ��a�A�ǂΉ̤T�H��<d�>ݖ���p�Ʈóy�%Q][K��YU��nQG��M6\��cb����vv�A�̅���w���.fI�E��|'a��jz�0��� ��cvV��~�_
��~t��E�|Ą�'1����(��$�����N%� ���y:��0�dZx'ٯ'�]ڜ�V���\*���彆�Pu���L��:#��v��޶�I�qw��ÀӢտ��*iQ}?K=Xw�8��k�k������4bv��b4��1ak?���(a�ۮ�xu7*Ǌb�|�4V<ۣ����:F��/��֦A �	v�{۝�'D$�I��ӓ5M\�IA�h�㸦��ooJ��]�[�D�*v��&ۡ�=���\��l5ZO��BI'
��i��4B\'�j�s��{�@F3�?���L�e�Ϯd��23t��"�
� L�椴��� ��A��Bi ��Zf��)1��ْ���׏᪞�Ri�K^D3ϳ:��]�s�Hȷ�KU�ʙ�M��9�õ���l���e\�J�C�^ �!��G�E΋�5^������u�>%�M1��KP��@����ڸ�A�%�~�V�
��A��`y�0��K_d�u�T��V�(��}�0>M
-'��0�Ջe�M�U҆��n��?�"�K���\�l���b�HY&T��%c��e(�HB����e����sG�}��3�m�T7���<�cɗ3���U�ʚ���_P6OW%p���
���Y��98']��d8�׭:bc3{R��6���B�ђ,J-_;�E����� O2c���6f��ʋz%ʔ{ޯfYSN��c �Mcg�6ň^��΀&�4��=_�2�>�E�o���� #��9��ˇ�@���e�����^鋴��k�ɘ��鉐Ye)`��h�YXO���f�1~�nN>ɕ��
�CA�Gs(P�Q�ED�1����)a���|8�Z2XWQ��5(f+I���ǻ4�e�<}���w�����b/w���8Uh�)��c*��98}-Ro��	J}a_��@0Գ!��.��z��P����%GAP_ik�C� Bx?�E�؜MI�k�R:�N'`�PnV�Z�/�K��+`u~���J�u/�ʛVu�@�V3������%u�5�U�IN�ۥ�Y��"����t�?ى\JC:�Q�S�/�9.��N�#
�U�S�ZT��S�V4��0�-M��2Bs&�i�Z޺Ce���0rJ�P� b�#��P�����^i���#��M�����pl�)LH-"�9����ka�����������O��qL,]H)`r�*:&��`cUf�%a6�a�@�<t�}	8"ugBB1�%L{��Qe5��M��LrUL���0���w{B I�qo�h�m�Ͷ���[|������{���̘-Քs�ln�a���M��c����J�ҚH.7&�?#���&2�5�M����]剡_ŉFzTD����>�,̀
5�t�Z��}ͣ�3 7m[���\�-���%z?w7��˻ʽ��\�ǲ^��ˍ�P�*��-ܓ���^/��6�I�,L�Q� �G:Ա��c�*J%5�@�2��̋�Հe�-�]ue�Z�-en�=��`mw�b�-����	�F\�����u�;k��\����;��cfuO����&���Ly�/LJ������ﴑ�����7��c��� '�n�&/_b���
P�q��cȷ7�ďh��yq�fx��h5��6���#�E��9�)x+ȡ��)Z@֡��]�?� Y��<�n�b�Dh����bA�>D�Pl�S�V�sq�\��b��p��4��{6ϼK�}��8�O3z��q�w�pbh�	[��u����Z�t��^A&fTzq�=;-����7Xi]�Lݸ���~��z���S]�U�Pڵ�f�1���bj���^���=r���k\n�t�����J&Y����#n�^z�ø��rx�k�7S5�	�A�>,v��zOѸHi�/��ٿ|����P/)�@Жn,\;��Ӿ�Mhx�BR���*�j>.���:Z�|EA{5�7<�h�����>$�[��;6�.�Y�����7Έ���vMG�Yu6ܒ����u|�qج]qZ���ݑV�-t�h��M
kȴ/�.��Y���J���b��Ў��4cF����q򫹻��_���}�n������%p_)�Q#b҇˚[�����Q0������8Ms�}����۔n�!���������4dV����8Fك�oϡg(G�H�)`� 1�t�L�	�%�]+t��&�G����l�rc�>���ig���l��n$�80��(}N���0z��2���e�IX4Kp��\�Q7,�K̗�n��L-T�����^=����!�_3���� �r}yGKl�v�lsx- zʣ�Z�`2�6����	�B��
c.��|E��$�N|�<��8��$P/�!&��"?�h��9l�#�p)FE7g5[��������A��D7����|9<�f_����� ���+�%�a1_C�L��\�Mǣw�?1ŷA�A-�ڀioK�?� �ҩ5۷㌨�%����j(��JE�d���u�Ҳq�M�D��L����}c=Ju#�8�P]�L��y�����.��1��P2�p��?O@#���{�A|e�n��B]to`���H�����舉},��/��%��>��:-߇�09o���r���>\�M����Dg�G��uJ��;'��Vla�7�b��H��"'�$�Ά3��\�����m�L�l����	eHt0��;ڋZ$��s��#d%��tѵ�&��8�:�z�Q1��O��E(O�����D��^6 �V��Wl�R�y�Ɵ��^M�^��ӦEaxH�s�+���_�V��˙���H���7r�B�b;�c��:*8�j!��� u�	�p �|�� �F}ہO�B�g���#D>BLh��w��N%4�K$
�?����E�ڿd���tl�\0]΋ �p�-V��ʘ�][L�?�қ�g�� ���1[e<�?	:u�S;�
O�VP�G{B%ܺ�Br9~O��W�8S�o�pW%��=��9o?�{�ؘQs4�zmt�����I׭��Uc��3ۭIc���T��J��LA��Q����Zi8+�+m��6{�-i�q�9oÌ�J'ͻ����hC_p�aJ�Qȿ],��q�&(�r�n�=vY�FԲ�a�gl#��'3N�"���X�tPXk�5��-.�8��&��D[�Q�(v�t����~�,�ų�D�I�M�N�d5���:5���Iñ��"��S�e�X�A	���_�0`���0և��m�������AW�A8% �)�E�/�L(��A��:䴺�w[Y/���?f���ͽ]�4mu�����B1��6F�!l;Z�)Oē�/��;w'�7�b�A����N0�b��{$5�\>��ON��g��|��.��Q��V���WlV�Q��(�פ����U��8����p���+[^d=�QW�y�Ti���rF$�t�HM� )̕Q���4z������i�Z�7�`��m#�s��~cV������]��`	�շ�R{6y �*����?�c�WH;\�ܽ�f�J̾��^��R�j�ma�щ��F��{L<��z�נ�i-G?fE�AN���َ�6��}��O��r+��7�w;8��(���m�n��ɡ'�$�i����%��1勵k���ak#�O���>� ��Xi��"o���A�++�/��85h����XspW�0`�t0����_��k���w
\�7�= ��J�ke��̀�^��P�]��h��{��D ��]��O��J�ߓ��۴����zʜ�����y;[�H[�U�3	\�����Ϭr�Ѩ�VEŎ����0��1K����L��8�(� ^���Xʐ�_V�1U�J�p9z+ױz��ܝڜ��q�����U��O2�M�QU�O����@Cʰ�G��L���^�%M!m{Yј�+��9FQ��q�y�$h�"[��%HGB�K���� !7�ygJ� ;�E�`	S�]�܍� yD)Շ�C��Nx;��(�C�S�t4�2JwQ��\���
���lw�[Ȟ:��&��zm��u������~
7��I�r�x���v��P��2b���xj���# ��i�5�?�ۅ�gѐ�XF�|������/u#�>��ܝB\�}\�x�aZC�kk؂_	�ѕ�'�K]b�0�����b�*J��q�4	�y%����Cv�y�
�=��	��5�-��QOnr�hjSY@�9�.#�|����3,ٞ� 
@���k]�NJ6h
ҝ $q!������X�۔�nv}�i��C��U0��u���=z>���'4����o�pcrw;�o�y�|����0 .�fDN�L�hE�P`o�<�"T6�]Ei���'u^����4l�dB#�}e�_��ۿ�W��x0[��dp�_�"⭐V-t�]�S,1) >�����jbw�6�Ü��Uc��|R#yH���&-^%���vQ"������`:K���Hַ�l<�I̿��%�$�xK����J�!���ܥ?^��_-k�>o4@6�@�Ń��`t�$x�˾\��uɒ�̈��J{=��
y�Y�9�4o�81�#�u}"˲�;�y�?����o�Aoj�����ӝ���✍���v"���s'4ȱ���u����q��[sK׎�n�'9��pL��[损T{~��N�|�ot̑�ͩ��Km�ƌ�����J��"s(�s�fN3���t&�_����GHI��Z^˧66�L�)CC��6��o�1���i��N�{�<�^v�-��ֽ�p
+���5R�z���
J5s%N�熂�Y�",�;9���T�[zq�ˏh��r�6���h�4/7�`<�� �l�P�dd7K�Eן��k^���˨v���j6w)͙��o�����S3&>��8�U(j���]�c�ӯ��q8ǘn��ai��A�~��z`:-���s�%E�\|U�@�Ţ���L���#pë��yL��ۑ��t���G O]#��t2:U�S[N&��/m�_�Fco�ܟVH�w�VKI]=*��k����M��+ƾ�fQ�tƺ4��F��Ŕ�����|�0�V���������>�dJs"+0k��xtn�n:�d,��O�'��i��:ç��SK�O�ۃ��u���K'�wHW�z��kP��+i�pXd˹��&S6^���Oӆ��6����ܵƏ2����s� },�;ܻHp���Q׌ea����-'� ^l[]�~w�G#kf3X�KU��VV����,��gW�uY��f��2��ɕ ��7�-�a��|c��U [�Ѫ�|,��ڙq�4��Md���C�?�͍Ɛ�j�|)aBD�� �E�2�ٞ_��uqN��۲��������q��Q�(v"�#�x<-:`��W����|$�/�+���c�Wu��Z�1�ȥ�%���+����	L�1ŗ����E�Y�,�f�ةL9II�#��������&�- ��"
(�tjV��bs�'�
�*<��ń#��ε�)b��������,I�w������, 1k������ޢ��[$��0u{"(f�	~�i<�����M橘2L4O`��JDǕp��5��1׮��.��.y8�!�o�[./���%0 l�be�yFn�_V���T����Z����Ph�xS��U�O���2�ll�Y��+X:Y��O&��uO�M>�iY�/�bX3�]2q����U�K��D!%�e��\���b��*L��AG`��gK� {�����L�z��!�G��Y���(�~�?�gX�Ŷ��T��;��ϙ�f�%S�N8�I^�m�x�u��<��+��O[WW'�fC����']�ܐt6�A���\�~:=��T�۱�cP��l �\	��J��,P� H�Fo��<�Eۓ7`�%�|}���Sc���ej����%��� ��Ɨ��4���.�M�SJ�dT�"U��M��������W�d��l���~�@^y�fR�n��n|��-F¾�Ch�ž9��Ĺ(I�`� ���������f$^_�B0�諮�o-z38�z�P�^g��\�\�`k�!��r��E)�/ �Tj�n�ҍwlI�� �Ճ�HC�T�?��۔��A,1�G��$������`��eY��	�n��+ٍ����R��A�$�\��-��������~��׏�l�:;�i]��33-�ۀg>/�"S���,�#+����[����
/^�?���{�]NMe"�ѹ�ZQ��L�>���Y���.+%��f�l�Q���6~���"Hh���؊`��;L��n^C:�s����ɚ��42gk�U��-}����H��(J��2��sK��
�w��P�R>�c�t/�>�M
�f��@:,�K��p�ʊy��8"��8v!��H]Y1�c!���W���7mpag��iao�@Fa�1��,T���𼿏���\gWG�	�0��n�湺��x��>�\Fg���'B>(�%'��=�,	s�˹�1���7:�a#!=gG_ž!,
(�kZ a�o+7��yyo��%̽�Г���`� c�SG� �	��j����y<��9!���'W'\�����@?�T��K�Q�ɸJL��m}?�V2�Ǧp�Z0<�:H��T��p�V8C��(�L-������;m�B�*��pꞇ�x>���U��� �y�ciɑ�P��ֆp]9ɵ~Q3yx�F��ǀթ/�x226[<�S�<�8�T*�ĂC*���eRm�ύNoCiF�Pv���2�d3��dK�kHEeL7��P��Ty1 "WШ��U����Ó��ę�)����X/��-t3���0�+J��]v?�B:��jb��Yl��B���K��}A��ջA��u���u��L�"2���bɟ��5����b�g/Jx����u�Y�1ڣ#�?B&�w�XP��D
�1�����%��<h�e���ʇ��~��Lr8���z�Is����c��R6��C�{#���Q���M��M'߳��SÐ����2��|�C��ő���zWm��]t$��/b���U��`\�w�X����<W��Mi�up���.�G�-HM�֝�a�?<�;'��Ï��;��pG9��T����H!("hۑ���7��c;�1ʝ٥�5>�R欤����:K&H�O'��&O�k)�?��ؤ�n���%���"��ȥՙ-�A㧴ێ��3׎��ְ�jv���G��<j*���I>>�i<|���|��x�Ӏ:#e�mn�ph|
���Ȁ���B���U�Дk�)�߼�G�����Q���a[��%�{����'Pm�:o��cy��X�
w�yz,�*P_��?=A��~;�t��Jc�&\b�hئ���(������e�:�T�S��'���T#F�� �dG:��\n`��k���g�9��ʳ���~o�e�A��a��~参{�ō0ȶ(���6��Y��/-�����O��S��1i+EH95w��v���F]��3��A�> �e�C[����OW�?�ur�����m#	�+C􌢒��[]���F���pR�x�U'l%���\��9<�G�x�Ӎd~� �E]��? �-�!3�L�����9����`h��qz��'-��ԅ�(�����7|bpf���ӼHz1��8�~5ѧuz�b"��u~N��D�Κtb�"��wꮩΤ�KKm�4�����kJ�0M�K �Z���F$��;���@/q��UK�]ܭ:�������uqL����}4��EdU���]V������fd%�H*��J���D=<>��{���f�է�*�r�|qV��(9Me>�o��=���JA��{�*(�κ�-�v�ӡ��g\��`*� l:��wZ�ZLt\��:U�Ǭ�y�yQC�����N�/��$���a�H6)������
M��fW�7��M��k�ƪ��J���6X�AqU��q`dL�Vv������ٲ� Tv���c�
�p�[2i����Sf�������40�V4Xз
����i	8��S�/:
l?�k�!��w�N0o;1D������ ��{ѼyS���9>����?�JSP�Fb ��&���TJ��K��TQDg�ʧ�B�8�!>�����U.T\g�N�}`&k..>�j��Z<a��m�.��r���8J>�X|$WT����æ�J��t�7����R�,��ȿ��=nN~s�/{>������_��t-���E�i��=���|I�y�$]�"�if���x��)Av]	l{�hi�;�k#��,���I��<ή�Ҙ�n���F>����}i��eI�?|�4��,e[�0tI����g(4�a�Ú���ݼ�v�3�';7�*o�l�˷���Ϊ�8�9�G%H
x+��dý&��fS�4tk\#|�!7��8�0����1/����^9��U��2���E�~�V�L.�a�gf�(?�5k�\����!�T����.��7�������D& U�
� ���`?Q!� ����(E:����.�����7!r�w����(�����������8��Tx�C��hG��<�v�$֎���xW#��z$�d�{��ǘ�2��"�E�F��W�L%�ݥ	����������:#r�Ў��nA����=B j�k������&���=�˿b�*� ��F��kW������2���'K�;�7�`DW��m��!+�e� $���g|��A*�������	1+��g��f h�A���m�7�`��BtZVJ�ȝ�u�Ɵ�U�-~ٓ�(?�H��נ،��JG�;]x~�ɢQs�`�u��
x�[�9�^q^��[�(fX8U����a_�헟!�eϤG��d�}�5�z�iLhLT�Oт��g2�m�㵞�/H�i�ƚ����N�^���A����M��c.ٶ��ϭt����	�a[��W�R�z�=S�����w�I
�vr���͚�V{Fm0�:��@*��8����j	I�cڞ�ɃZ?�$�C�I�������f� ���ɼ�P�l׺�W�C,� �Y+�O�I�,���������Ւ:���/�'4�A ��^L ��/���T0G&F��"5���}�z7*y%Od{Θ �ׇv0��>}�ձ����<���]�T̆�w��z��6���߶��Tty  U�ܗD)��JӠ�P�0�Mk �7B�W��4`��3���W�3<?:��x����6�����YN����s.��&(��ia�Q|�frn�t檖J�܍j��z�<�Q,�ڥ#�4(>��'��0a��K����pao�� 	��vo[��%��h*��� �ew� ��A���5�(�e�\`�|g�}N�l�yZٔ�]�'7�#��wJ-�����:�]�V؊W��|Q����4��b�����T۝�7�R��!sF�u���S��.:���M�Hϴ��[sH[�bbel�"�|b���AVTa�v��W:�C�F^�cK��C�;я�E�P<w��.���':���ᦱ�if;���ǋ�Gah��9P
�����2��S(�53��>UT�-�ΛGЁ�F�ޑ�8?��g�'^s�5�M$����,\?���`�m0��Xr�ɢc&?�� �Q�I����������FE�tY�Q�8�����X$���G���4�'��a�5�(�ym4�5�tw�ȡ/_�&[.�1shK�O.�l��{y(e���\I�Qt{��A��TT&��%J��"�R��Ο7X�Q�����0�%QSB�J�U�#�+܅j�,��_���wU�B�{�EJ���+��Nb'W�Vot]3�4�
�\�����S��=�g~��|����=��SʫuZ�0O�{�e������o`�@�E�7�o���d�e�l��\�}�@�?��*�N8���u����b<�nrr�����q'�ˮ?4��_��G-�/�� �)�_��=&"ǔ�QM��u0�%�T����epP�vȿ%M%�ͨ��$��Ǎ���dZ�>��T9�kXdY����N7f��V+Bj��r��N#2ܻ�v���E��uBP�h�����u��
��?���	��i�|J��8,�7ݧ�C�P���c �o�� ��k��k��R�cDm
Z�[RY/�OML��ke�U���}���
��w3�꫊���e��Q@*�Һ��aL ;j�u����'��̞~��Sm�r�>��9��2&��S0��2�b�7��<�m�����{�>7=u?@�v�xJh�샱�s+��p!��Ѡk[��!^��5��V�L��&�h�����m'�ͬbS���'����.�}
y����&%�lv��2CC���ަ���m	J������3>]:�dR��D��������'�vQe�����E���R����}M�_�b^L�rB�ZIA�#3ֈ3�(��Y�9�gؘ��!cc:90�[{,�#�&�.�V[�O���0�o}���a)Lȭ�1���1��)�����/���6rH�H'�,�|\�Y6T'a�$��9b��P�9��e�,r
�}3����`����Co0NU��h���(��!�"_�w4���|�}��(�_�>���/KJ�x=#����)���[��=Hc�K綌��~A��?ɯJ�]���-�d;������X��]��AD�V��ƫ�D%X�����H>f���e%JE�J����6�z�SE���$�����ij�}������]-��!�w�l�RLҼǚ�eC�أ,��B��R,�-�~>��s�J�D�9�d���~��NW�r�n��lWwV����hכ9hmp����C���c�6QٯO��c|�Ʈ^<��74Ux�m�s�ߟ�-7n�;\t���ٗ�D�O/�[%�@�o[�	!��Px�5*��Q��G���y��$Ӗ�A��MG�K��9(!�CM����A��&��O}��-"�����>-׹C�1[B�"��fض�ݣNh�ԿpxS
;�k�����wRq��[���P�a�V|?�n<|���DsUr�XV���Ѭ�C����)�@J��c�C�������o	9Z�>�����
�hx����x�o��4L��:-B:�S���ÕA���\������z��k�%�s�8!���x�����2��_ n�x�s���Z(V96��N�@j�8��2x�%=�&سL^�""2���	9x*��f��%cB��X��1ն���T�b��o}Ea�=����o�e#�(\��/4B�#wH	���
�ּL�yL�LֻN���/��x1ـ9�u�
Ƀ��kv��~��:���F�D���p�j��ό����-�F���Q)E����%вX"&�Kd��F&(�I0��<�`���*�M�������p�cT׃���ʝӟ����@/3�ΏsÎWd������h���W��o\`��¼m�h�#P��Ƀ=��H��h0;R=Շ�x�����x��l����6�F�Reѩ\�-�]��T!�4�&읰|�4���5!/��}yxp��SŵP����&;�6�nW�qg������S��E����sn���SZ�'t��FDh�[2*x��R
k��Pk׏�r��U+���?;%A��\�6	#�iQ�����3��΄Y7g�|�{v}`��DԨ.x�4F�������D�	�g�7�̮�'rE�������_=��(\bx��(N�KAq͖��?�c�U�O�������ӡ3�}p���L�V낽��"�.���;]/�'O��MC��ls9�ۈ��/�ִ�Q�9,	�4Ub�5jb�(��={3�D"g(ԃ��, 52�Tͯ��P3�S�R�`]`�y�qړ�)��8��<��xc�����W٥'*t*F��vc`�	(�/�^�£ef�Z�%E_PП~YCTg ����b��+ۮ;�X_zW�ł>kLO�πdPr����O.�&ႀ��yd)�t���d�W�"I�14����F7DUS2�����v�OE*{�����F0��0!������(
��N�S�M����)�??H��-�k��_@�w��\X��ș!�4:�1��'�Z�)X�>�0-�h�z�|��2)½��C@��}��j�
�Pr9�b��H�2oT�l�.��߬����ä/�QY��h!���O!�pU�j�r�|  ��Kmhx�H��
V�&ʢ�D���;'ڡ�u��\D�x��X}Lqr��0b�f�"j���� M_�V}�%br��pw��%Ѭ��XȐ�	e�����mBt£��v+�Pz�4�s]����vܓ���DDu˹�߲m�w]�O���b�̗�@�Y�-��^~E�-�D�$�APlƭBSu��n�}�����z�MJ�o:]4	x@N!%�L_F���hl.�y	Ai���l�_��l��1�u �O�1�9&uj눘n����<�e18o��k�b�����3^M68�!��ii�����dǌ��E7�h���ָ"��m�q�I��:�Ɠ<V��2Ư��&h��Ϋ�f"�.�M�=�aЪ� ������CTµ������u=qõ�ٳ�;�БX�XW����������> �	'���F��i���Ϝ����&s��`b%���-���NZ�7 �����͛>v7�<��G�L:LV�o�/����C8C�s�9�eSB�)�)�to%;������g�Wn�U�<_ �����N1�
�{���!%�]�?��2��Z3/�$��1 ]rRw��E<��j��,�!uK9�Z�K�A��;:��_t����N��]���d�ˍ�+�y�Y�z��!Le+���ZLr��0|� !��uxE?M\\�ֻyT��϶�Dt0���5���R�@,���rb;~�V��Z\��B��7��82��=.���_ZA��O\�Ig�<*c���&�Hn���P�f�� ��M�E�x��X=Pm�L;�!��4�!0'EC�$εcMcM&(�E�u���i�i�p����յф�v�)k&�(�c�90�U*O�K��t�<.��������$��㳌�H�򽌢5:>�:�I���L�pX-�tw^���������7��I/���[ro���1��]O�a�T�K��T�'`����_ٞ&`Y�|�W;T�7��xP� �̎AeUd�}i������.��l7�Ow�s�dA���_Q�X]����������c�����-Gȫ��W��O�,���so��w#��Fz;* V�7D�M��VR��� �cT�l�B���q�y�%�DGĽN����`0P�Whv�1���缮���׿L(�w;����t�e���CM��𺄼��!��K��lQU��4�Jd����-A�[a��B�y8P�TDFe���Jc"��׸������&�S�
<�D'�n/���No���w�����`IO�6��B��w�����F_\��H�J�9�����K�z��-ׂa�z|z����3��Bc�������u]�M��R��Z-��#pM�1��}�#�PU�5a�YE�~$�,%-z����R��N�z�5�Ǿr��~���#��Gۍ��7��v�!�.֪e�����Q��o����C��퇓�9g	�mk?ь�,����N7Qs=�~c?wAq�'�J��Q#�7��\+���P0�*��V9�����qQTÚy����t>t�U�si��;���cꬁn��葷7ebq]���>C~m4�0.��l�/I�)��H�!F�>������g���P!wH]K��U���ȏ@����KO�#;�RbΌ�/�[�+�bϠ;��|�i��t�Aph̑{�,l����'��)�X����1S�	�S�b�m#�����������<��{ien;��|�AU�@qd��#��ѱ\�"z)�����������W]`��Z��k�U���`��G�4�;ٸ�ν�Ӥ 1�~�SRZ�>���G繞�2ᙾg�@�=A7�x���[*�'0�, �N���B�1X�A�;9|��<���BT��a6�\S�p-���\�������L�2����v7�΁��;�A�)�M3�b`.V�<b���*w"�5
��sE[U��(�������`#vy<�m�p@�&�������BO1]꧈�c��r���ѧ��M���$��`��1h/f�x��-����YP.�	���fOaLʌ7���F�+�z_��.\���p����QA�W�Y�׈���Ƒ�A����P6�U�h�0�=@�uH���]`�\�ݢd��Ĕ� ���wa-_��@�.%�[�xH�$Eͣ*hŹC{�8^6�/�5���	����S6�ȝ}B�7�HFC`/�F[��=2��q�8��J��؄#��? ��P�e�zDH��<���H��ڛ̉ǐKN�وj��k�8�)�Z�o�b��FMj0�m+� Q����+��BR8֛.y0��Ѿ%Py�c�2Y�&ѪxοW�QS�S��?��r��c�?�b���m7��@le�	�ё�{�W�J{��t�-����	��~�|t<�>����.�rV�Wm~/]Z����b����m����0���6��#w�*0� ����㑗���]fce��&���y�82m�=�6��(��/�ճ��?�����l�ࣿ�2��ǉ(),B�(�ɹ%, q�{�"A��+'��y����@p
��	�e����ZOVI�U'���*zz�c���Y��3WS��ږ$*�e7���$%,"���6�fFa�*S��kK:ߕR��Ӷ|��:Ȅ�@�ps�>� R�	Ĵ�B����G�P������b���ܽ�/�knk �NYO�<+��1͑Ek^� o�0}�B�e-v�E9�gx{��q�>)����"���_n�a��I睙���`�F�����A�e��O���-��AUY��V�5%h'1J����Q�H3��ޒ��X��;]#<p>~�G���)k�� ��#��w��ꌧ7�ʔ�ӛ�}0�8J���r�����H�9$,�b�/������e��=�1�+ {Z	r��{@H��X[�ٖ�M`������r5ު�Q�P�S�R�\�	E|v⨞X�g@������0],���%��6,9���$�>BT�mo$5�IF���/��~K3XA��H�w��O7�P"hD�b�-<�u]����K��Y��Ρet8�� �_e�|o��,;��§�K8]��~���o�����^��H(W��S�p�c�p�~2Z~Х�JɮT�:!${?�G����j��9��2�����c2X�׳ܧX�k8�辐�!�4�\��U��޾+Uf�_���H�H6��x�iձP�J���b̠69s"IY�ů������O�*���[�oj�-8}�.p*�����M�}��e���<Σ�T
Lc"�R��a���
ӈ����(�M3�Wg�>6��L�VɈ�Apըdkȟ.��19(v��Q|Fh���V��.m�j���V�`�7	pяI&*�v�B��˽0g�nw�=BR��ANg�i~�w<�����kmځO�^�盛����C/�ʧi�����·9�N,��Nh#闝d28u	S���l�{�T{������ 5�0y�?[�΄��x2�J^E9��n9(f�3�1���҅;�����P&���Φ-�-s^(��,�^�-*��S�jQ�ԁ���\y��T{o>xG�	?�8@Jt����������������bULC����z�!��9ٟn����kG��!��Y<݇�/! �|��w��7H�J.�Y&79����>� ���g�{\���7�Mi2����0���Z��G�$���~�A���<���4�o8��b�g9:��@��l
g!j�Q�#���7��f6�9���i�2�N|��u��n�3�.���ۇZ���3]̪_q��cM1��`	[Y�h��W�qn�B��!����Dkd��()p�
A��S֊�OUyL�G[}m:�>�rn�*�c|%|�w�$����[k�T^,l�i-x#@%=co�s�iUN0���x*���
�S�`5���JȪr��`F�z���W��x���d@��`�����w��3Px�R���wC�MCm|���.�7a=�G�7|�f���7�juT�6��ne�&߁�Eաx�D��4Qb��0;g�о<�[@�F��%h�P��M0���CO��U���N��z���|N��]��lAhp��xG�J�3��S���p��R��L0��;�yޱ�������8P��ө���{�6����z͉Z��$xD4|��#�����2,	���3%b�1�p��q1^b���ScW(�^�^Q,y4La��`P���F���وݸ��y�l�<���q@����ו<j�-�V�p�1K�8�U\�ŻWN�-�����e	u��cdEo�S
߅����M@v:�}-�_�b�O��"c��嫁���Z�������Z�f�{���/6)	T����(72'�@d֑F�n���wN2��r���('���}��Q@v��ű��!��+n�W8V��	�x'@d�ʅ?���'lV�����Z�/�m��c:6�LP,�$kR;T5Ȗ]��Np<(^v�9k|@Z��n��Cإ�K�T+��K�b���w3��JrQ��.瘈�	/�H�|Nz���x���i��ˡ�va�Q:ʆ�����c8F�Kҍ���g��K�ReS�Ş�3	x���W�[iXGϳ��z]j}p�ҊV������sM ��zD>I�L��9�JyR^�홾�]k��~�[!	Nr�A�I:�-��roT3��5j�f�� �
������I�5�oA��̂|��f���{�6���̹[3$��Ɏؘ2��m��'�.26����|�����`�+�e{�N\��1�)'�n�����G/#�u�ҏ(��>[:>G~�z K����4�|�n.S��`��U�
8���ڋ�AQ����33�{c9��M��2�3���N��J��@�+,���-#��~�l��]zsY�ْ�*�Q�A����Q*�*(�Y�3h�*&(H%�y�\F�:/��w�_D���cj�ߧWD�(! ��o�jf�@����[�"���ց'W� �����vѣH���o�� 6N'i.@Y5���1�����ś&�
��C�L�'�L�/E7���"F7���d�T&!�9X���QI�����Y��6/NK� ��\Ѷ7*7P.�}��Y$#\PP�*!^K��a<0�)X��N��e���1v/�f[BYI��l`����E��S���/�B�yB�Fx�� ��DzX�>�Q��Dǋ�Yk�|싀%q��kf�4k�T:����	:�c�m��X�S۾'��C;�	�S��*2��ڞ��p��u���n�Qt�Rm|��*���0QL�?W�C��ݖfr�&Ԉ�#Y�	_y��˪Lę�*3i��%���c��UX���PM���U��k��>�?"&�9a>���{�@	�\�#S���x���_ʯ�r[X �}���~)�4V{�m���}]�k=��O1�ϞZQ��M5�qQ;뢫���й, ��v�wS���	�y���~�w9>�G�a���WBT��'/�E�:�K��:��j~}[_�o��u��ōt��{���>hR,Y[s/��ÝDZn�k�4#,R�
wɳAN>:��0�~_��)� �hO�������=�i%d1����L�>R ��w�*<;u^�RcdC!z�YL�R�9#������w�^�#y������r�zd�-埓��<�d�͠����I)�V�R�d��U;���q*ߐ���7=�.��Lz{K�=��E��TdCn�sh]7k����Vbڟ rgC�����Е����n��B�Ŗ�E�`�2ء���"W���~=�9�9�����YLA_�s����|�$�3�2a��ؒG�^L���ԤŹ���U\xZ�β�{��2����p��2f���$�o�<���Z�^6/�{dG� "��I,�Gߛr�q���f��Z����G����P�����Q���$��<[m��J9��OZu���t`��;?-��52��*��e����7�:��ū��������KFN��T���\�&�}�MVQ���=�ݏ O�)l0*�t����&�#8@H�s���g��z]�r/�0Up)$�2��h	a�J�3�Ư���F2鍺�·�/�@=B�#U�u,�j=\] �葇D�rryͷ�w�X@�4�O�(��v�i���.*7��"0i`��$+�ĕmrR�z|.|G䠺�M�&5�ڒ�K���7=[�c�>�{�*"(w�Ⅴ�}���9D������D�-��J �#�|�Gr�PD���:�X�%_IB@�����Q�󨥅��?�!c��2N�IL���r�1�m�w���3�9����2d��c�c��n�����A�bcmV�K�=�W�$̧_#����r�Bw]Br����d.��3�RìX�u@�ha�#ܴ�U�^-V��P�FU�	Ϸ4�|̭�Ҵj�> �5 (.#�!!$�Rn�n�,#(�����z����f;�H����x� �C�N��Ħg%�⟝r�VZ$5nӘʔ�,�,�V�����n��� dU�E��⤈ٸK�~��%�6���T��r�>�Ar�@�1Nh^ۿ�A��?����; �6�v�ǉE�K�;��4�%�g97�fiaĆ!��v�Q�%S\��L���9�*7B��+ҜN8)�n���eA��}�RK���ާx��<�"^o �6:v�<��O����(�����L� �$8�no`�LYr#J�	�~.)��ab�r_��)tD����#x�&���Tr>���F��t�M���Y����։��6z�T�K��Ea�2��S}Tv����`�Z�7F���ϓi�Et�?�����ڍe2���Cl��7�r}ig����g9-I��*���b��«�t�[(X�K�i�)n�7����0���Zߥ�(i�S��ޟ���y��nr����$��=P�������&���Д��γ��\���ziX��eYȃ���+�[r�Ͷ!v>t�ҡ&�ۀ�S|?�'�gH-2=�^ZP�0>�291��^\�+�z8+��p��Tv�Ws�4�P^?��)��b��!x��0����C>�i<@���K �7+v�F?p�D�4�#��EE�1Ū�����j��+�S�G[��a��7A~)�Of[���� Cq1l�m�x~�8���c��2�q��T�mޠ"���)����t�9u-6ҁ{��7&[_/3�$�-|�;���L��M[��g� ��e���݊�Ld�O���J��.ÅO�I����6��Y�\hM� 
�g_�1,�t|�����P.�%�0 |U�����R�h~����y��M�r�����݋��Di����e�*�ۍ��P�5�yp���)�UY�u����-���a��s���t�Yʌ����B�7�
����y���%�v���j9�!��oOw��F���aU�ja�
R ��.��	�<�o�j�ٯ<�}�k.�L�B�vr�����%�&�>�p0�5r���*ϡX��E�E��(m'oI�h������ۢ�g��Y�C�g^�ʦ��9{�f՝z��»[�U��	����>��p)�z�n�.	�<��\�la��� ���X����fj:���$Ϣ�̬\5/Uh]k�ӽ=�1t��0�-Hr��wwz!����w���u���I.h5&���i�Л4V�c���h�d@,��R�sJ�C�.�}��ϳ��,?�w�q=p;b�&���-�.���6�e�W�cĖ���V&��Ze�
)�.liɹ�F�[��N�*�K��g���D��$��V��	d�(w���[�;���&W:�\t��r� ���!)�ѩ�ɐ��B�D������c��M�ː>X�^X\nB6�/�a��J�Pi\�~ڈ@��#:�4�?��=#�#�xŔL���Շ���,�jUY���H!Õ	��\�;b��{`/>f,Ƅʉ�΋���\4�0�jm��iˡ,���rq��_�2��	��4�+"�y�׭�-���*y�C��i��oP��Ay���ȭ����'{�siRhO%�d҄��̻� u�Xn��w ��B�������\���b���o7P�#<�?�I>���!�NN�*`��>/J
 ^
�Ҿ����;���c�4 �U/uhY��&�v�½��4`��Q�,�i�q�,	�iV
��}5$Z���|��-4�r0��L��ƌ==�H0����hT �Î��V��4ֻ2��7���$?���6�)��)�:,��}��G˞�&!�D�F�����j���K3�eoB�3�PfQ���!T�y��4�?�m��yr�E���5��z�ws�?�B�~t�o�����_�P����>�z���$�e����/�x��m��G�b�M5��BǊ����;#�-��ݴn�4�jv��G�� �fr"4�'����b����qDXw/0���!W��w�r� Δ=Cs�L��瘘�������ŋ�rX���nv�B���r�s��{ݺL5eX��{�1w��A��/KyY�	�ى�@���˛h���]��K���Y���`��U��)�a�Z�¯�l�}1�6�G��2"�W�N�2���nr?+��}�w�Έ�w����[:���d�f&o�7E!���!<�Sʹ��`�ZNq׳�����V`3�P�ۜ�*v.����*:59��/Ch��ؚ�I�-|��[Ä��k	4�,�:�4t�fEǤ>[�[�����z��vZ�����m~HO�pi[&l��$��Ի�H�S86s�	�E6]��6+�'�_r�>ux�j��|=?πp'����_��*#��=��I<�o��)A����%�&)�+%C��}3�-1��K�Ҙ���b��Ǒ�c�wZ�KX�u1ڶ�y���n�wx�d�oT��=�����|�Iq�6y��d�e�'~�I�*2��$h�أi�cИ�}Vdi�	WÑ�,Pfo��!H*T�4��l9�1*�\n�|��PD����ծ���ۓ[��0L~�+��:9�@N�s��^n0��G�_~�����W��0��6��OR��y�N�.�q�$M(Z톷���,r1f�JIg,~b���S'2�g����5�����/.��|Ұq��x�*�b��i�^�W��MbZs1�i��b��c���X��|��&��.-��y�;�S��ᯄ�d<�ʽ��G��oJ���G���͆=	���dE���1s�F�!7��D�x[Un>t �ip�6UF��^�K�JR�]u���Gde2V�@�ҳ	q��S3b�L��S��C=Y�b�Yb�Ml1�ܨ*}�Th�elun���K�0�?���ߞ��n�W5DV�~"!7��~�*v����#���=�`�=���a'��+�@��"2��b1��b$��\�*�P0�
������a���-�]|92��2����q���TR�L:���.,#v7�"a��Đl�O�*�شb���W���ԮJ���)	[�%��T���PQ؂qH�`޳Y��G�Í����`��!@!�M�N�G�ø�X*Duv𬪰�s�q����#?���&��}� �S5��ɾ5�)�0��'	�%�����l֐S=�7������=�_�.+~1��}Q]����%��P nٮM{���^�Q���#�} 6�zLH�)��.�-Z��d0W�챟�%j�zڋ�ٌ6M�����	HX�aGvJ*\k���ku	�23��w1Dz��qy�3@�k�L��'�8˪T	���;+r�,��o@�@$s5]�n���x,@,��#��f��{�E�)k�>��UGh[8�f1�A^�xAm��%��5�G	�#qF��UI@'lj"a5Iz����x@�^|�R�/jO���l1�T�~X�r�rA>�� �_��Q-�G���eo�f��<A���
�z`��?�/H蝨��!�,�ưA=��SG����|�CpK�9~8-�
k�	_*���dl��U��C}���Ԯo��5�*�^ԉ(t֣!�X�&�z�L�8��;�����I��_�-�:�W�NF��� ��N91c�O�NOxgt)k�^��K�L�}�N;�p� ���ƺ��o�kၯ��;a��M�
_3x�Y���W`|�Ę��Q{�m��6pG�9��8x�Wf��8S�E���a�Ł��U�l$�`�X�(���q������>���������~�q��D�*�WO^��Ɨ�M�aύ�������,���8j>)�w	G)�������t�ĩWZ�_�K�U�D�`ʂ�-ᆮiP:�����'k<զ�*�8�n/sA�+o�4�Ɣ��WX\F�z9�4,����i���y k8J��y�
~��$���fr��fK�N5���3�2I�l�@���8��ԫ5e����J{�<}1j�`�o�"f؝�q��UG�C�

b���."�	�����L�z�s(cȨ�85|���;��P�o�E֕��������C����&���m9xZ� �l��uYtu���\T�+ݗ�J��!�X(e3oE���AE Q�k��F��8U"�ӭ��w�oU��:%����?(FB��TV�m�)�K͒/��	.GM�l�iWM�3O:nWфzRA�;����I�s}����KXx�$�~��a*��j�s���\���t�I�;{8r�#M]*Q���&�55gdhPaY����]�{՟F+4TL$�XD�t>�,z�Mդ�
�W�s9�!�0-@Q�Db=��(�� �Ț�mv����ݤ�
tJ�O��F��u�����>�p�1<d$ş�ᣝ	*�������I+��"٠��y?���Tm(���`I�x�2G����RF��-�&vI��:����}?87�W��2x`x������	�����F�z6����d�Z+YL>���Bj5�H��5��&�-
�
w,��ڕ#�
V�x4�NRm�[�kQ���m$�"2�a�s�ןnAnl���%!\�.�����Ip#�ʗ�4�� vm��h	��x�~�y�J��!�X��!&6{�v�8;�q&�<U"j�'�E^Ŗ^�mc�F�=��{�8�]�
�@X\c����'����Ε�J}`�B�g/�&̚����;���+Z�5�����5���$����4�"O%�N��Bf�y/>w�w_�D�6�b83l������"�c��m���l���2(T�V2w�����K��_0��םB��������Y�)��եq����*���6��P7<W�3$;>��6���(��]���Zi ��%�����rilː�i��dL�0�� ܠ��+j�q�.��;��;}`A�m��5�#X#y�QB�P��(�)ϰ�1���@�z��Zt~f�c��G�&t��:��G�wE��VSK;�	��d�iG&3��Z�z�P-L�W7�g:��d4�v�{M5��蚫���0�;Sԣ�t�@jX���q(�iL/�ͱF��
?f؏�o:�5-RB�e�"�Z~��\��2ܸ�bX���Ӫ�V�?~7��nc�O�\�*'3}�l���'5�f�ى&G"{��
/#�􉹈�����-pm��Sy�2�>�#w��L�W�HD�TO������x����Z�&����]��&?]��[��������������8����6+c��|��TN^�I�}`~�o'!�2nUf�_�k�
��\�)��'��J��+�N��v�T��q��o����h��a����h<_X����TT JCF{L�Su�ɏ2��M&wyp�W2�/Ps��S��V�!����X���<z./�P^���so���VE��Ķ4�ɇ���t�9��_IQoH�֮h�0x�	��ư���i[e'��-m'x-
EPD�j!������X���63d_�w{���T=&�+g<�f�~{�;n��Y;Ӄ L��=f�����tUw&Km���̬��)� ӥ
�c���wFUD����{����ˆK��r�b�:c����
�蘢�j�wK?��
u� ���W��~0tc�9	��%�3������Mlq��k�x}�Q.]J���^Z�[v���
ϖ��?O��RkO��9�"����]:/�٥���2��ᘗ�E���b!�i��(pG�93��I2�l�B��{50����iGќM=S�'�&����rrY|x��m�rf�ڭCj�f���~�;�U�Q���1*��wO�y�FŸ˔c{5�h_
�z�Mx����@�����c_�T�%~��Z*G�
x��M����6���=�ム}n� ����]z	m;�La�;eA�߆��������I�`-�RB+������`
�,��;�#��g�I�Ę �>�O^ϱ����s���$�8~f?T`�����D�ҫ���`��(>\��� i\Q�d���(�J)i�4�u�U�;��fk�,(�O���>����J��֚� }4"Z�j�D'b~�?{jyj��L��;�ٿ4 ���xGAݟn\��q�ٙaT�A���f�G�� �Y#�C��Cӄ}��N�s˸�9�)q7C$=���; JP�Ţq*��i�j�-�$G�e���#���RA�/-��eN�v������/6������̩|��ߊ�w��jW�	-�m&���1c�T{�23	#��7C�%v��E�h�ñ�9��;K+����_̞΋��b20o�e�,�[%�c{��Ƒ%��6�<�j~���:��;!����'f�:�|7�?��U�26pcrKw:s3���$7`��\ȎSj�����i��jG���R�Z�-�vp/X�q���%?\csv|#�PQVoe~���#}���Uh`��}A��Ǔ;��q���X�u�/��Ǵ`�x�t
�g�9(oU�r����\o^������jU������`�V�Y�5�KTȊ�e��0���tK� ���#%��c�iB� ^�C�g���3�I�"�\��T���'�<WM]���8K�H?"��z�>��W��bC�(�#pW�^�/�i J �~هis���6���E��r��˻�"+�i��%~�6V�:ըj1E�����T� ѡ/��XE42��0P����V�j�z1sW;p��e�1z9Br!�*����e	�o�g�g�/�@fr�^CMv����NPu����!p�|��mf*-0'��^?���b�O��M�Y�L��k��蠳�Db��f��7 G�:��R`�b:�M�2
�� ���v$�*����s�0:K$%���)��2��� p��E��Ϲ���e�th{
��O�AV�Q�O&h���'i�1��̡�禱�3�CQ����؂�.E��H_� T�l���Y-�$؋��a\�� |�\}�QI� ���W��{�d
��]�8��z�죢�<��1��j̀��Q��oT�d
�?EQ�7�(*�-�e��������f0I�X�F4ѳ;7����(�r���Q�^'���}�ȣ��.=��%C)�Z�j��W����o�������,�s�ڤ�駱��
���t�W,D����j�۰»c,qk҈=,���/@M��́ә��W����qIٰ�J��,�@��e��V�smh���)˂�F\���=�����f*�R��.���Xn#�2�H��wd�}Yv@;��	�a4��
�a;j�2,�դ�@�jS�#�Ch�+&�#��6���/�%�[�����]@S���%^֬{$��oN��c+�zÒIr��h��#����B�Aty�d�[�2g��'812�N�v]������)�V��DX�U�!��a%���;�
�~�~�eEF�I�+w�"h�y�X���#+�;T�S(-��E8)8){�W����P#�U�P�b t�'0 E�[�V���`1B���{c�'�������"/�"��㈍�:AZY��(��-&B����@#�s��]���
�W�>�O؏��ª�XmL[s����{I��e�vmoa ��z��]�c����ǂ�����m���4��m�Ǉ����l����E�K�6����9��&���о�vI���
�z�\>����Ù��c�%cxݴ��(r��o�����p���������Iƒ�>��f2ϖ�eñ��~���a5�&!n��,�E��F��x����bM�;-�!>��_�]�SXZ]��*K�Z6s���CKa���=�~l�؅D�����9<y����/��".���P"���q�'�V�o��e�C0�>��]9�\"�l�b���N�[��)g|,!x�~p�hl��0Y[�%���ۉުӐ���V�Xm.	jѵ�N�]���9�s���@]'��Z�U�D�X�p����z�Sѓ�`��"�Nd_����SX��Ϗ�I>�hriG��L����c�Ĕ�C6�����	���F�� �weD��Ē�'�{>��{��m�U_�ʨ-�zM�C{�!c&L�q�گT·G���� �툠���zS����S+D���[�>]��[C	���~n��*�)�]^���	���FC�ù�M]na��A����	v�K<V��zf���ȈRsŢ����-�;kC�v�Hj���Eoe!hp�"��D>�Ҷ�ʂ&��JD� ��M����<�|���p�J����l���[�"���-<To!��/�d���3W�O�sm�͝�gw?��&��߾��}��z�OES��iIv��o]��f���jY믏��Lx'D�8��;\�bFv�28
=ͬ��,`%��Kd�
�1��:�̃QE����O{���b6g�㍵Np!RѤ�!����G�x���mY�G>S:�)8D6gmI&��2��T�&%s�\T���Oz�?�t8�QG��̕e�ge�)I��a$7n�z�3$��@�M�̿NɣG�e����w�s\"j0�f���@W���.[��^q.���G���8��":�ѹ��g���-ârں��@6]��U��M�M��~�6]��e0��gƷ�]C|!g%�h/d��#\������o��qR(qI�#�:W:=���#�{�Ӑ��!x_���čN�K��=���9hC��q�O&��d�OB�g9N��Htx�T׍�v�3�z�^������ iK��!~��r3�Ւ~C�q��%u6
ןc%��R��{�I�1<�{#7kDr F2�*�c[����T�/��{�M!��(�Dz/�\�~��B�(�̟�D��
�U��%��&�W��y�Z$'~��� �M�
�W�pF����{��'��OH�e�q*Nlu�6v_��%\�W\@`x��c>+��bX(2���kn�@{�8y7Y(�"��-�,|�ʅ��d�L�#��v�(W���]��9�fG��]�T�?ݖ*.��X���Ds/vL
��1��'w���lEF���ZNb	����C�؍󷖞l���% ���uFu�_�
�m�L Q�t�Q���s&��ʄ���ӕ�}�Z��
<R�Ɵ�~���I$/ݔ�y�4V���{��P��"S"�0���`L�&�zRHYՀx��N6� ��6�˕
m����>�4h�=�(�8�dsV�ò!��oc�O�
�����f�����O����dReNƦ_�����"ygC�a5Y�\
�;z`�༡+�?���A��H���_��L��G�pLO�䜵�-W����[��� �>U�*�"�ZoKK�Wi�J�C�=�n�b ���K�d��,�y�F܀àv����j�jBvӝ����fŦ����$3��v�R.�J��=��Z+��e<Tw"1>�ґEDyw���4�w���\	U�F9Ⱦ�q�E|�Q�&���׺���Z�e�74�pV9ԟ03iљ�SŲ�QT>g���#�U�1!�Gu��̗�!�n��W��LB��gu���H���s[�jo��B�|���ҴgY��)�"��q���R�*P$J:�N��P|�{@p���ͷ�� e���l%�?CC����$�(�6���L��/���d����i��?J�Jz�j|�5��Y�����l�n�|�o)+��/���I��Q�K�J�'ӜG�L}����Y��	��Oh�0����@�����x��e8��0 �w3T������g�DW�Y�g_R��T�����Cz��e�r���v+E�99y��J��M�e%݁E���B��ĭ�D�J5�Q`�4 �UI�j{8�>)xw����k	�������=��6��u������@Ʉ�7�H/2F�L��\1lW��M{ #W&�Z�nż�)�y�A'�!�f� �v�Z���/�<���Y~K�OQEZ�HÔ���0��V�x[�CmI���\ �7dX�'7��8��m�h};a�[cl��2����[��W��Q�M�[yǉ'�xs��`��!�@�-�$(��*pd��`����^���n�<\�`��U�ӟr�%_}�T�̵�W�ar��f�_m'��e�M��
.J�W~
�{Z>&�t�Sr̎��zC@l�o�Kdb7�o���<h���Ak�S��ʈ`��L�萤͂�p��N=�������?��G��t}lB}�j!�Yfa@�ϵ@B�c�� ��B
ca:�� ���W�-�� �ù@��ƙ��=L+�s�L������1��1�s��qǅ��  I�I �z$v��U �,"�AL���ĭ���L��BCH0G:�Aؼ��^�#?���z���	x5xOhp�'.�Az�H��� =F!s�7�o3����f�h<����4�%����{l���0� W"t���z0�ģ���cw]�<��~��~��No=����΅Oѫf,��H-���?�E�B钸C�Z���M�y���b�3b.������㩾�]KL��q�B؈��w����8j-��ܰ�{[7�aqȼ麃��~4K�n}Wvi�L��<�(a窥�������� |(�FД���!?�g�ǰ�w�th�M���c� �W�-�쇲{Y߈�n�v9<�
\�r�E��*D_�ꨚ�e-ږm|�Ȏ�S��7a�^d�iO�i����%O��>�����1��]	�T�68H���XY���l�.���֏�2�Zo���1�59�!�۳N�S���^������n���'����<G�l{�ۈxf���F�1�=�c�� �mV��-�A��"���;�
',c��<I�Ёl�x-�kD��������j�j|�w�5��(/#W�O(���}s��-z8��X�[���E*	* ��P�ꃁ�i
����{���+!l�A��o����ɑ���Ȅ�r����3]���eاa��</�Z���0�x{�c����P���b�ij@�Y�F91kB�ǁ���̕�x���r<?s�b{�0AZ�,��bU�s X�򢖀�Y�eͼe�ny_�AAR�=*��Av{2�g	i��p^I($�j��<$� k�rߝ^�_%�������"�'$�_`��%��P�w��� ��s��V������ �G<{��� j15e�g�2F�T�����\�P���r�\�G1�x^b��R�Ό�+������ĥ`��#p-��"@iP�]�0���}.��=ѦV^9�=X|�L��y��]�*f2��G	�<����j%�#���@V�"8�׼�u����ez��R%n���n�Q*�ۮ))�E]���~�u�*í1�0�X�U?�}ғ(c��I�U�Mї�շAϣ��k�x����tg˴%�b�m7���Xf�+�n+ۖ(r��ߛ��W�/��/�_m�BE�Ih?Y끭Ԣ�헨IhD�=�k�ڦRM��6�~3�3vUT�D����el���B*���E��'>hS��1:T/�'L27�	zb.�op.�Q9md⬨��C-��J��8��/9�(g��-'�i�~w�� ��͢�P��^	d\X�f���[s{�W#�>��G��8�9CD���l��"n�7s�0��(�~��oV�/����3$�~�"?���P/�]NЄ��1�'�	N)��x�aS�f��c�믊b����'U��٨��*x�	T$����2�
�[�X�Տ{�|MlGUiJ���V\���l����Asb}U:�)	���Vb���
�눎�x9l�B%z�7hPK��,N�?�%����z7��EEk���Sp wP@�`v�dOz�~7Q��O�ˮӕ��	\u�vY�˩�C6<N���ߗ�s)F��pE�Ѻ�Z���ǳ�/�l�D�ߒtF������Ӳ�k5�o�{h���Zo�"eW�Z���
�%��J1;5��x�閻P��t2P�PU��ʹ2���@��4��	���Fa*VK���^�������$��̀N��Δ$�ڞ�H���<L���k8ՒJ:s�	!�s����L���5�i�!�=����"�����t9���./L�a�fC��=�U��'4��OYn^ ���|cK���O"E��D�O��h5]R�ş��@!ݢL�nƵ"x@��Gnw �`��eY3x8��t)�k���0�ͣ#m�&������ppX� �hh)J��ھY[�0�zok���[�~HW=��r`@��k�Dj�KV-L���\A�;�<�Q��Ho"w��,���e��-�j;GEá�$p��[�_b��������MO��1�{m�y~�5��^��@:�8�v�e�燊	u�I�Qo���ri�'»d�1�s�����t r!�!Lq1���&�I���5P�4M�XkEg2�Ru8M������o�Y��v�M�+�N�KU������R�R���=Va�<��-v
7�^龒t��r���),�闒C��/�z���nu�^�ئ��!q�Q���2CcR!ݻ��Pؐ��+C,���t�{P/R�c��:#��Z:1sO=�՚�7��񐫻h���c�99�/D18'
:VO��eg��Y? D�Y�x\��1�r¤�[L�e���ܽ���o�0O�\�l:��h��K��c�g���Q:��.�z,_3l�q���һ�g���d�I�(�����Arw@�Hǈ����]UZ�U�Ri�e�_d1G]Kz��~5DBu�$(ɚ����lA&5�@�^h�l�8v~_x-�S���-p#��� W�����������e�TJ`���\�I�:��aЀ����	��iS���D�UR�� �b��U��?_7q϶�������\-6">O���^�H�K�ܠm��*�����$P�m\�ҵ�Sk�]s)ƕ�#�8�����ܭ�ڿ� 2?UI�6�/�ݚ�>e�2�����W-�P�6��/W��-Ӫ(;�l�ó(�B�m��L�0����/Z"�@��hO��@���6���|��l�������/�ܟD�|��o�z���/EdB><��ۜ`}ːhGӠ��:*��qՇ'�B{�c }A���q\cͰSA�`�?φ�EP0\���9jz��Gy0��	��u��Lg0��2�⴨!s��l]kM����(�̗���\�{��wqW9��O�.��~���<N���Xݲ���ś'�Eᇞ!*&DaA�R��D��/��Ie�������"yv�����
u��R�Af �~vm��[�}Օf>��v�$_�
��W򃊷ٯq�r -r�y�i'w5��/�U�i���HOl1����k��]�NS�x����k���^H+�R�++�do�}q�k&>�=ğ�;��Ř�Сt��*�27	q|;.*ѐ<�؎�p=�Q��u}]�}oͪ�y�����@9�`n=U
���V��6�
�(�1aH���.U�r`#)��CV�lZ-��m�������=��W�b|/���T]��'m�7�G�'=�u�;�S�;N�KPe ����OU���JG�y:@|§�������TJ�mk:�� d~�Slx"� ��E�fW>�?!^�*�{_)�N#bO�zфg�+��D�"r�+s;��}�C���U*���sW�u8f���L�R�U-�s~Nөd`�X:GQH|:L̳�k���4詁���tѧ�b�b���R\�l��vb�lt%�cW���6>�v��Qj�u�ėd�N�ct�Ӓ���}���#k��9?	�+�΅s� �5�.�V�B�E�������h����ږM��p�$����z�~SYV�� \.��#����l�4�9�>�����=,�iT�Cԃ}z8�����t:���c��*�x�,H�##��KXg�?
l	�h9W߆���H����&�:蘛�w��_��U���Y���=r��	]�{��Q�;�y:CʭX�o�2���N����~]2�1�	��H��i ���|%�)=a*�p�����5׆h�#=S9��s	�ȳA�����>ݕ�~-~PW'h1[~������wЋN�������.��!���C}�}p4n�V��d��V���q�w5�		�e���)�Ρ`��(�7���ή����G ׃ ����~.�	�W�#�l]!+cHog�8��#�W�f��~��4~��yU; 	U�Yo��ЇHT�	T+�t��v@Ι����3�vZ𣉁��,�����<�Á�t�ڱ�C���o�x~�=��C6��"
t�{>�,�5	`f����=?�;������a~�7����1�B�`��ks�I�K�l�Nk���u�$ �2��Q���bנ�����x���Ѭ�7��+F9��M��qA	W����5(`�}~����Ow��/*�3ڜ��&Ge��`7Z�ރ(�4�FO�M��'Ds��!l�x���Jg ]Qb$A������A�d���x��1-:��6}�HЍ���vgY헥��a�\�|�m�YI��Z�%�:E�>��D�3�����|�>����mFw��g�U�K��B^Lh����/��a��^X�h�����,�V��"���=�9�4!�C����H�����N�i�"n��̓�����W,/�Z�ܳ/�@=WE z ,�c4KO�J��#�gaŵ�==_������[I��E��~<p�B��p
�[Pr��U����4�I����a��Z���lW�v8rb0�z+�G��&Y� C���YL�m�XG-Z�3k���W���7$�`�M��6�k��F�	����qhWd�U$舻o��n�D����ը��
">�޽�ՀR����y��f���ŹTm���7(k�ٯ���#��~�*�\��e�xu��^�xj��́*E�;���!�G/��G更���]�2��`�A�ׂv��J1��.�f�b]Z���Z���T�%Zd�BO'FQ��ϣs���� ϒ6�4�ˠ�/2�I�kl2��&M0��Ul%f�7�A&���\g6����V��؂xX~Ǆ���W0��ϐ�2��ؐ��GZ�a�!C*汪J7S�0Ņ�';� m�X/��T|奿U�m�WX&��e[��Z��WC8�Z���4_�	��Q�C(��<1�$n����k�2಼�u;��a��=���[���p� �V̇7�bZ�2TNP]�q�!�
A?iL��#w�"�.k6r~ᙢ����3 }�'&�L�K!l���1P�tv�� C��U�k�~��<�N���F�Yo�e#�����"3����`�x�̲V�MO��f��o��$6|A|zr�&��CvJ[=�7\VC��[<�n���N��9����q*c������{/Ȃ�&�2��/`ρO���ޚ�V�`��w�6�3���~](11	�BZ T���||���+T��N֚�i�z���y����I�G��i��d]ݛ��w1 �[��8&x3-A����4���1 ��%Uo]�o�T��0���L֘W�T��nV���}�`&|�3�!��V�;b\��N����'Xmuf�Y�T���	w�=k��?/A��W����3���`� ��5|�*5΄������wb���5�r/(�''	{\���z:�v��� VA���g���� �4cu�������&�Fv�e�k7w�: �R��;k�Q�-���&�"壺�"-��E��Y'_|D�L/=�nl������� �<���./�rÌ��en�q�y�[l�?ނW!� �V%�K sM����>��4k{B4 ��b��-R.<)�ΗPoF&h$G��^?�%�"�"h�#����w]Inջ���mm$�	�K5�դ�S�[���r�����Z�����=�V�0��nD7�0���;��J�[b�����7#���[j`����jB����bpɻlD��vx��N9g9:=�L[�$��V8�=(!��j�}�p,����U�A��E��� ��T�!�Ey?�v('T���r�򰣒ˀ�d�"ޒ��Ȕ�� �.�ipl!��ආ��,�o�<᳏ݿg�8�S]/7.��h�*�����z������������5�ɒ�wC���� �Qͨ
���{���w'�r�rF
�Kc@�x�������G$��F�
e! �'��J�J�4X���}U�L�����&�-a�Q��3���7���w`_CV�Ĉ齞�d�O)M��@�Dh����5T��d�<�e��Q�!!g6��ɝj�I�H
p���;;�l>�e(� ��E��{�  �jO6T�tz���Jѥ���*&�2:��c���e��:��~��R��26��X
����O��:����fu��s>C?�Cs]�xA�R�F4osP�\�	a��*�b� O��Gi	ԓJˌCeۆ�o~����45��{�>?
�"�iٺ�I�|���F-���g�u���A̹2v�r<�����Fh�*A_�����_>F]���"�+C8a'=��I�K�W)En��i�K��qR#L��+���wJ�Q�8�9rT���j)���w���yy�zE/-z�;̼$������.W]�Y������b5f�#!�	F�~�+���TH�{�?0��ʳWxS����t�}��m�	H��tH!��zq�Mi��P�������H�� %M9�;�7�	�R]yI\e�;?��^,�
��*rwc"��Gi^�E8K
f��Ov�:q��V��B,�Z������r^�� �G3+�X�y((�vEcc�j���3�q�����i9w��-$��@4[����xN��P�%�����{�jޖ`4O/6e�-b,%�!#�h2Ȑk�ط�����/a��Hz��0A�?)�'�M�p������a�h7��{�"Ԟ�^c(u��q����<���J��ڦӐ16+�����P���p5N �)�p@�]?�7L�RKb������ﺥ(��_3�*-�AxUkI�krZKD�$͇�m
�~uH~�봅����/��s�8���%)w2'�99�h��k��_ ��_���;cgcA,����}�kO��uT�-n��2Я+v�0��S��E�'Q��s��W?1�X5L�/�P����������k���d`��P���D���-�������*3HC�L��]o��^TG�'�O��s�#|�3qXL̽`���d�g����6��Э������`�7P������϶2녀{I6������H����]���`����~1�t���4u	O�e��S:��:.�(��Vw�ۥW �b�twr�ܩ���iC'�Ӆ���^��ΉZ���ٚ�T�����b�[�B�K�E�w�"kc.�+�0�ja'�ﮖ�S�]��_�����yH��t_�	���_���Ll�Bz�s�ˑ��]����^T˰��I6I�#oR�ς&g��ﳝ���\���|�`��o���2>�[v�����3t��ЛW��';� s�*=��}\�1,��uh�AC>D9{�Y�	�)���3Nˏ��Y�ǅ+_ж���a/���y�3�Txt�1i`l#�+�B_ܒ~���`�)'��;�(�Ր5����	�/�j/Na�����:o�\>Q�IDf�3��w���(
�Rl�Z�<���C�ɛ�A���x18�|��(�ʐ�p�1����O������ՖpS�=]�-A�c�O����<���6r�S%=g���iC���d��z��	[��ᑸW؄NÐg	fU���-��#)��p�~��l�B�o�@�4�S�{+�{N��_EۀJ�FY���Y�E�H�2R��=�a���}��.D���^��@�7@Lo�W�FIF�4�w���b�h��j�M��G� {��k�̆߶"D<)sF����e�{7J��K ��ު�L�s(���A�� �吃�{S��{ ��*�TG�6���΢�r�?ѽK԰���>�P�*,�Ƙ�p�W
�_�3|�"g�	c����Ba/&U['���p9n���CKي^�t��a+�8V�x�"&&�f�Xm0�5X�l�Z.o��Ǻ��5Nf+�/x��`�ajY���H��N�����&��`�MvlC
��	�t������� ����1��o-\�ܕ�ˋ��;��p}Eoޕ���0�D�ɽgA>즡�A��7�Z,EZ�v��5
�R��D��r9�lC�ns�
&�i㎉T9�+ <���aI"�6��yeO�ٚ�p��O����#;����-�Y1U���[u�:�=�k�9+�SC>�z�z�x��H�W�)���QHe�F�K�����˃%,��F�������,�S��X?�WHݾ}37 �zZ�X	���6�a��\[qk�8þ0�~?���� ���>�jr�沼| ui�1%��>:��?����3)m���B�ߧ�a�~�Wx�&��?Q��]βD�Q��9E����H0}����FP��8	�3�6���2![����7���f�J �׾]�(i�'�\�6
F�YS�q?rLF^t��b:Bj�?�H��6�Z}ۈ��N%1����XT0��Хʹ��;������_b.��ơ�-e\���9����ZL��R�����q>P�6�Ӌ�AC���0� .3��(���g��5�I����^�� �������S�ݷ�f)G6CU��� ������}��)23yQ/��Gg<��Wq�V֍a��˻���K�tAGg�-R����Grn�3�8�Jڦ�U�mQ��9���EQh͹���_ke<�����V�=�'�) �:J�uv/-6uɰF�m
K��vmM���c�M5l���A � �M{�/���5���!�9��,�Q�#J9�+�!(�s�)Ǎǥ�;���&�d�>��r
�N��؇�/\о���j:;�L�rQ���AjR�S���Y3mxUBA���g����b�[,�:���L��nZ���7��P�7pd�/E%�Oh۵^�Ep�V�߆�U hiq
�'g;��"w�qy�g>|���SjK%ʄTJ�3.]+�b���T<Ҳ?�
r���N�6oH���䦽���`-{J�D;먦�����xk�=���^�{�=2l�KH6���1�i����2�v�^vq�i����Ox�
�����)O��A�t|��܉��e��'�7�B���[g�Γw�*��״&!�\)o\-��yuv�}J�?���DЕ�J��s��/M�P��k4�qq~��`�esX�C|��A���c/��k��c3p�����S�L�@+�몑 &b�4c��5Bz�H���z��I���e``���W�#Yܿ	I8��̕��tzSt��#���8�e�@��m0cXY0� ��5��D������r�lBL�E��U)RC��,r[u����K&7եv���|���my˧���q������9�^1+���Vo��ثQ�
زw���꠫�8�I�XRU(�X<^���+��Z���>B�Ig�ϳ^gm����M�$>������U��6���<�̼�Q]:����;�\�\m ��1{n@ꪇZOPd�n��6��
QvF�c�ɂ><�� �a���*6�A96���x�踰G���B��8��z%�^�Y�˼o��S�3�0�n�/D����S4���p�r�Ϝ��̜�������(c���O�МП7r�.��4h��u|��ig>�J���׳����֬
��3�ݔ�w�D7�K�'�A�����3E 7ዽ1m���{���V�<�~h_�-�����=���ک<�u�6`N��B��Z|�4-^�fc:h�ð��r��\��@��@�-��Ҝ��5��h`�����o�~)��5HZ���ʔz��P0!��t��7�]��U+Xo9m��E��������qOv�(�~}���S,��[}M�kY<F����{�BB᱔��@&���tI���XԽ�*+��P4�P��LfE�D_�A�Z�3�Ӽ�ѵ�f�c�JC[
��9n���s^�v��ގ�˾�z�UXp�|���Q=8i����H��^��S�~R����N����d���۴J����h�F�A7���H���晳W�z~c?v�_۬��u�D9l��w�ޖܨ���D?
�t$D��cɏF�ag���1��M�
���˪~���e��9�.��ѓ�"�=��/�"yRC��.��3ء���~�>"��_�"�����:��p9sv6)��a{s�Q����^ag`ѱ7`|�N��V
��)�ү�cz�k�Pm��`���X�T&k0�� s 45;���Jx� 0
�4%4җ�cA�S�֝��^��yn�W���jO+��2A5���Q@X! �
�+���&#�c�����qܮ�̫]����w��{��*M2#��FUR7\캽�_Nh�rL�^�Te3���)�VTLDi +�z��q<R�+1������0Ǥt��4�R�FC��Z>����s|Y�7�C��%d~�u2.E���^vn�0B�0��4f�����Y��kM������9쁴�:T.������ygL?��¥��s٠rl�IW�Ȧ��,��j�N5���[��3�}��6V��o�uU7-��Y��E:$6�/^�|�r���+�1��N>�C���Gw�s3'���&�cn��ǜe��O�c��9K�\����i���F�Q��V@%Z�����n�1Wr����v����7(�K�a[�;��q;�:��n��P���ud�s��9��1Ѭ�d��蟿��X���c�)U�a~�kL�f��dxv��=�\;gX0X�`�H���()W�K	��h*H��o����Fwm�S*�W`���'�>-��	"�(��&�Z,5���k����-Է�ą����"˷9����1[ ��=�����rHBU#���m��6 ��m�_���D�)m�n}�!A��^_�64��5i�Ȉ+W�7��{uB��� ��Z^�il�I����zwTVi�� �#�]�G��5�����i�	θ��/n>_:����w�VHp��������g�Я`o�
v�m�s���H �-�8'3MO�ACr��X�$�J��^u����%t����U����>�J�`�����O[�E
'`#P��i	�Er
��U�m��F���P=i���U�(�t�%.8G
�y��7+"������
��d)=�O&�f?�2'��;'�>h��h�A�OݿK_`#�����BT'Q��n5����eSgol"�|�"B�sϼ�:��<Q���e��Hd�ō-�܃`��:���lx� �ο�hωJ����->g{���R����N�ԩV,<\��_&9�9&���F��S��rٱ,��뫕�@x��ӿ��痏#�7#��7�mй�]�ebj�i���3qR�y�)�p��:��诗i_*	:��h:�@ĀU�~���?S�N��)z=�ˡ��K<�"E��+ꅌEw6�LR_�Iz�l��|O,I�>��7���nE&���' �I���l����5]ӧ�e�z�����2��mtw��T�<���~�����h�|�sMݶE�=	M�Q�����ki}��μН.0��B����A�np�A��2�L!��q3BRD�+����O�n ��7��fХ�U�G<;���s���e�s-�_Ʌ�kpb0�1���9.V:���ۑ��X�}�4'BP3�I��'�7�lwCn.�z��d\7.���v8i+S����6�����4.�X�J��ŜZ̚�A�:�������x`E�Q�ўL$��ll�&�����ٲ��`puv}7	��[X����B32a��z�>]Gve�Ʃ�őViYP-d*О$��.�Rh��ѳ��(`���Z��Y9ݙԦ�mqT���� 7���^��]�Mm�o�� �o��ڎ���i#�.+������i�-픿]���,�WM����熏q���ƭ�'ɞ��2�򧫗}�jbη߹_E)�z$'�w��x�&�GF/$T���F���0G|����,�21�P� Dw'b��'Vc��Z4��x�˚qխ�#�X��I�y�`��<ԋ[�f5����Ԍ���u뽚�d��zR��������iA�WNA���ƴ����h�O�=\����r ����(W/�G~�Z6�2O~���t����mKV��AQ���'_7)1Y0>�����kt4�/���g�8�����H��A4�b���(����F_�0���W?����ѹS�0+���U���Q�: 5�g?��p�P���m_�mb{�w��bCuh��of'�~�sI��/�Fs!`�ӯ0�T\e�e�����}�@x��V�Y�����($<�dI��R�[< ��K��{t6O�I.v�[��oys�r2O�{��όz��ђMx�[�������}h��)���^����-	m��+�A������x�`?͓������J��Ɋ[�!M*�5ń����D櫄y-3k���DV[n�*��.g!D\�S�m���UC1a��L�s(���ۤ:qT~;�j���}��FuO��`%��Ʊ�,�)��Q�G���t��`7�>�%?q����l%�7X�������H�lo�ۛxc/�ݡ �&�>5<z��j���z��^�^8vq>nE� �fb��9�UefQa��,]<E�}��ݎazzǷ�q�7hG���!J0�g�X�`
�[��>ň�Pƃ4����u���k9b橭�� ��t-bB�YğQ�.Em���}�K*���g4��h�s@̳�����ԣ��QF9���;�9&����0f�2�v ��u�����3��q�&���R6g"���K`�M��C#��bn����9�*�HG�Fkđ��Ȱ+M��L���L�Et��l����k�E�0:9�$���	*]���J/'�k�h���sM��*�v��Cw�F����\�VI-~{з zg͟�B�![Ob;��vN��d>}�J�$L	����:p[��7�b'��/���f�Ys�[D���?�E�AX�tl��Jdw�� ���Ǝ2�����MTUaT�(�O­�ٳ�q5D��?���1�Ӽ�g`14���+H�Y���P��3C���Ѧ�+��Fי�W���O�L�J�t���l�GMYL�_p�>�5L�<��\Ѭ�ۭ��1��ц����t1���5<Y�Kŝ+׺�:B���,9�J|�Dd�a���7p_mT��J�a�G�jT�5��9�L�p 4"���
y��L��T�	CZqQ^@�'�l(`����
�v���^��I��iw> ��[,l�Y�)�����v��D�H}aK5ܚ;��A\�]4ະ���ڠgF����z�I�&�UQ�.���]C�dg~+�b����ˈT=RQS�¼�QZ�Y�Ym����y�,��K������^�­���� ՒV��g�	����/�e�s���������h$Ϳπ�W|8wd�D[�J6���d�)�$��E��|s��x�#�O�r� ��������?�@�C���W<�����7zA�k�6�Q��FgHeeI�B�����n�P�4��Q��W���������zW�8��?D��q rk��Ԛ�g����>z��n �Oٻ�� ��Q#~M0!���	���U�S(��M}
_Hhs�Um��a�I.x�j�[S�U��Ci��s����p"�=�Qks8�2�h��ڂxt��y����z%��!�B@����t�Oˌ�I+��L$��r��CFO�V���R���wc\#�i�Zy����n�\��h��ٹ����������n9�<�[>�Ez#�w��%r�]��)KG(���u���$c"'>�q��p��{��}�=���;.��Zҋ�ovo��z���1�:�C#k�ߟ�Ь���}D%�㹉e�ڮ�#24I��&��2�*p�����f�旸�r�l�ہ���ќ�������e������q�56��WR	-]�7�c����=��wa�eC����Y�aZ+��!�$4/[t��SfhT�度�n
M�0)XH~X��$}�8)���/�?B_�<HY�X��_;+>��t��#��x?����%v�׮rF�Z����0�
N�M�2�~�Q/���T�RPH������~�!��U�TG)1�-��a�[�Ȍ���oc=O��~b���Zw3�L�'|-��x��G�8�t�p�OiC��//*7��1�,�G����b<����3~��Qƥ��>a7Ύ:���$y&x��K�d)G�㷏lYin
ϙ���M$��lQc�툈9u����2雖�uO�^���&���y����)ߌzԝ�9k)2����"��<�<JW�/g�͞�2E�疙Y,j���LE�e�h�n̆m�sO�vS���0L�
��7��~�,,>��a	��Tz�'�u�T��.�#ߪ�������|vN�B�Do�ۀ�̅�2���ܶͥa�7�K�`dt������'@��0j?.�$l�:�]$Z����Y�ݷ��7,���QhY�Há�̟�'3`{�^q�~S>�(���ba��+�,!�!�K��k�dE{*�� Rs�k���
Z���H�8 �T��p�W���N�d�����V�Y|HK��tc�|��_:Na�{��E��K���bG��9C�_쯖�����9��� 1�B�2^�y���M=�ތ�����M]�R?�n�Jl��wS��8|�".gX�km�*ܨP���K~�+��Ԯg0�_���)L���
��^�{i�E��n���ڛ�k���B��bl~6��˯7�Jk���d0>��ի�0܂hH�"�eX�t�VSE:dBbeZ����l~�.?#�˔��I��8��Cݸ~A�1`�y�E�Ɇ�Η��h�_��M���*�g� ������O�%<_ѓom79��<aO0���F&�ySu*��*
?M���>��-�/�h���Ļ�wg������,�#�S7��)�����ג��z�<�yO��	�i;:u~PHz߂ =M�hs��DM�49���)4Ӡ}d�ǣ��/w�a��!�[�Ǘ����!�Wtwd�]%��Heu��m��E-,�i'��f��9�5�)0�ج$@�@-�`9��h�gH�|�}뾷��(G+�DC��Y}QJޕ��JC� .�a�#�8��U��_���a�Z ��~l����N2V�3�E^��9�^���HJ7Y������Ӓ�Y����Fe����*���T��6a��|Y�lwa
�:�p]�m�i�$���$T }��r�����~0_$ X�F�_V֔$�\�����_2�0���MIv�v�H��a�wC#���_�3ėă͏�C��1���2J�?�4�g��Ǘ�%W��\�<�C�a�6E�hn��m�%�ZD,M���w�|�B���mm&��8��x|
m����O��=D��D���eħ%�V����Ezk��Z��ߣi��Σ���y�s��ëf�0K������D�J��� ���a��R�2�C��p���Ą�P	����WqR��e���&h!���~�"t�w��C���*^R�	�JjX��|G��T.n���M*fJ���E��mV&�Ơ|�l�õ+�:`�L� �Tm�MX�=M�g�,�*+~��pr�8:\9����à��r���R-R�MH!k�(�O�2�L������}�g�~h�Oc����tkw�>H�NG��dnjă)$i�&p�C(
����29���]b��3�Da���}k��^#�8�j�{�����m��CvD2��g�gi$��©?�,�ڵ��z��l����[
�J��v����h�1�Y��j���~�kP6�^ɯ٪��B'e)���_ϧe^"F�r����l�h�� '�8S	�2���M����a�Y�>��<;B��?��Djئ�叓x!f+y����~�\�w���ƛ�hq6"Tk���`��n��_�&`l��ã
��@�U_�i?�_���h��YE��Z�
�Re�U����ד�^��@vo����Ή���]�"qE��a�J�Vy8��tU3/Q�Z�E�;O�����
��;��|��K�a�!G"�^+�'5��l�!Ŵ*�YFu78��p��a����<��6_� Z�I�'�iAW�}�)�3�fpF�e��������ՙ�������X�wq��_L��0���4]�f��^w
s� �q�q��Uy!���9J����"*"Lר�6CFբ�G>��D��S�q4�1�UG��.#�"�]>ɸ�;k�����^�G��>�$��	 -�&V�Bj&K贂�S�:�7��\�N㿹�$1�ņG���/��A��&p�:Ut6�YV��a�Mgh��EM�Xrq�#�"$&�Jy������Ww�����c�:�@a�_����&�G���ф�A���a�>L�!��Z�VN�s1A�;�ɝ���3�}v:jP|�I�(�	�$E����Y�|jEb]=P-7����P�Yz�M�(n�������ѥtӚq2, Vy!'<P�"��y��{L��4"�#�L�ā��0c@m�qI2���F�&�K I��YIA�W��(Qa�B&�p]7�_r�$A�()�W����ﳅ; �9����t�
#�C���vN�S�O�N�]\��r��� !7tbs�&Y�K�5jOG��2)�,���;�Y�~8�k�N񂴝1����9�WO�S0����Y�[�U$S%����XW���Ȕ����+Z�Վ
6۴{�D����ْ�����C�&�g?�ْa1�a�Qզ��4�S����%vm�B�<B�(��?R8�:ye���Z+���s���������������?.�ф�~���V�Cs{���h�;��$�HW�W(�Xn�L�b{~��ZI9ZU/��j�u#�
z�m����`�vB��>n�P(�ܜ��0�n=E?$~2l��#0���m8����5n@�$>��=y�=�p9�1��^5�ѡ�-�y�qw��B����O�x��h���\~��,�j���f�6O?�d��N2So���>'y�D2�f%6Z�MƵ�`ho�bV#�Õe�c���w���Hzh�;^��_���r�2���3M��t䀝���{����Z�����)��3��Q��"�%���)5����Ux����_P�A�	��ը�/E����N<T��w��:�|��'�6w6H����2��O�����u��c��6M��5iEo$�AG� ��JB9g������pzU�Wuƴ`-��+N7��.J3����
p�@	z��ON�:ZUc`�9�s3:p��?��4%�L�5�&�t��� ?۩Ηc~�d9��~[�X��i\T��G��̭a�e�*@N�x���G ���z�#ڍ����d̦�4�7p6��F@l$!la�Q`v%(����
�_f�WtM/��}tM*b@�Z ��2��uy`uQ��E�:꽁ȾV�у���!��}*&���Z��5!�z��ܥ�W�e�?�3.�/����#{�?`N��-�ə��!���(a&���Rٰ���ۖ�Ъ. _땈Qr�8��H�H�N7=�R�*�5!fs/��{�'�t,b�v����Z����l���1����X��Z©�w��/�F���f���0���c��Ո"�xa|�xw ��=_�Wl5 a�ainiPR!Y�#��d�&������0P%��$����vE}�^��G�-��������E%���=Zk�%s�����8 �)�Fi�W��h�B�F������plpth�W�!�ia�V���٬vJDqȳ��
��<��2�/�È��9D^pؗ5��u(�e���Ts)���t��xEj���ʂ_�U=��ic� ٜ3'��)�ݫ�;��,��r֦�;ip��7�KE�Q��=>&@�SOܫ;y�r`ו�kaLa��R\�`.]e�J}� ���
�����%2�����;n!����zqc�EM����"��|����'�M�(ˣ��W�:E��t��%��
.��V��f���K ��

�����"��rU��p�G��d��Au��0Zָ6?.���VlNM�������#�$ٞ
�c���??��g";K���#�d���e�t�!ԋ���8�JT��`�$�.���$
Z����WE��"�/���	0���`�#f
>�ъ�yE@�*iXHzk����eM��������#�2�*�iX�#�@�)g��;`}�S⢅/���C�1�S�K1�s�O�j��a��Fq��ϭ�\B%�,gQ�D��n4������-&��y��nk�y��\�4�sri�֊����N�v �q�mOZ9]J�a�	�L�?���T��q"Hk�K~���;-��Y�����_�
���aY�"8&TBv薬�zp��	/� �xY^��'�b�I��nR��{����"���ؗ�b��.�nԋ�!��=�����H��'����|ՁPl�d�ҕa=є��a;���5]Pa���e�y���x�h�=b�1�[��Ǹx}g|I�+|���W�\l|��R�C�$�|tD�V�8<�arX�"����O�H�_��C�z�����`t��F��s��k)���˓��4�U���M�9L<e_R���ȹ�뎿|�����}W����<�pqB};����0�R2~睚	;�݂$<d�&M�K�	�RK,�����_��f�J
��a�K��^K72m؜\)�}8��:K���Ń����:���������o�� h� Z��S��T6�{�Y�5��F�T�U�&n3����n�l��sˬ~�f36���ey�V=�=de�G�^-�*�1�5:������a�Y��M���t�mTU�+U�̷�����&f�E�Q�V����r.��|�:35��(ː��b��(��n�?[��Po�O�]�֔< 9rC��L��d�O����pB[����aa�(g�o�SB�*_:�������Z�k���М��y�p��N���@{��؈C`G)���Q�������@]�S>2q�ˑ�6�UJ���/SGɅi��v��ŉ��n�k�����#GN�LR�B��з����G��m��R�^5 &�g��{㬦�!�����+��ū�� G"��!�&��M���:ԳhSa�Mb�k�Φ��B5�I ��Q<�/�͠#v�����0|�@S)�}���5E��q��6�>L+c��;���gC:���u���F��$��jڊ�BMg-k���t�E۶� 梐v�<�$�����b������v�-p���)}��{�}ZE�?\tW:e@jk�����A0ٚ�ݾ�R+ݟl��O�<��M' ڶw�\��]�߭փ���Zo ��ǹ%���j:��gu��K��ͥ$�p�v_1nn���Lx���8K8P  �$��ا��L#�oUd8����S$�y��?ajO��
��]�ap�Td������^$l��6b ��	��?2L�5x�K���F]�)e^�Tro[���x����v�̆B��\ƬB(���06S�HQYQR���-�s��b-� 	�&Y@ڲ����\c!�<�1�qx7�@��X�8�2βn�Ɖ+qP��W�%o�����"хNQ���$0�Av��r(��X�{��ȶS.
��XD�֔�e�ف�9���h�o��c_��y���!5�_���/9����i��;�o��|�/а�����3����+�d/����1��B�wd�;ɠRW7��N�ӣp���ʹYF�#�D
�y���S�}���U��u����z��@���b����'3�-KAo����1-γ�b����[~i��b��J���Pd�fr�j��=����N��ԟ8&r�"u�~���~����F�m�?�c�t�ք�Gy�VҜI$8�U>��k��)���`�a�����]�/��6i���{0X�A���f��-�� tm]CY��(�F���Y�F�ƥ���L���}�Z�d�te�Uer.�U��s�xŤ�0��{U;Ta�{[���UÖ��(:M��J5+����#s���a�ވ�f�:�6He������uwѳQ���0<�.�i@l��qVvp���G>k�X��#�6^LK'~el��y�nC���2%��a��dE��iS�yy�0e���<\��*�%���#v�#Z�c}<U�籬H���>�z�Vl��[�V:����v�Q��s��xP�qb����S���Gʑ�cʵp[�K\WO���of���q�V�lIw~�_f�U��nUC'��fwTk�:�1E�sp ���0u�eԝaw��#�Pm��UUj�o��j�!��󊛅�LXC���4�g"L��:I·e����|��OY�-��'�Hw6�0�B��D5���6I��^�y�!/ݲ6�9~�ݐ�����!
�6bBG+�hbu��`��<S��V<���_kzy���䈭p�� -M�,M�X�P!�������L
�����i��)RXl~jR�)��ʣK6�f�\�xh��K�r�~���F`����mdzca�����U�|bλ��(�4��J&��_��1v������_���t��9SL0�+'I�ā1(���˳�x����*%Wլ��U��5��*���?��Ķ�y [	�>�P�J�yC��F��QU�.�1�X��(�<��s4��]���F�w�����Ȫ���=��PPQs?����A6� �,Ь�PN+p����j��j��5�I��[Ii��{��xJDA����V}g��F���&bSX�#�ԙ���N�$�Y<
��+�#|dp<��w~A󹸍
��М��ɝ �:�C�0�Ě��>����ϔ}E<�v{`�c:E�m���?�����~c,u��NE�mf���]����YR��S��;�C�)RuM�B�T�[�f~;T /�0�|}�����њJ�Y���,<�M��F� �qY<�F�����!)l$������7�J�ތ�.�G�����n�]U�O�~6�@)��71#l�q��a���.+Uw�Ģ��g��aM�>"�I&=���j�. 3ϧ3�|��=��+E�U��w���d���yVHTқ��+2�J���(x3��?�,#}���h�X,	|�zKIL��8����f�Sp���Jd68	�� ͋er6�%O�_Q;cP�kfp��k�9���w�p��<{F<�#H��蔸�26Ҭ��b T!fn")���ux�@�*ȶγ3�c�5~,ʞJЩ��m��̺��5L���-b( Y�zA��WH��׼z(J#�[����s�����>_�-�J]��؛�l����/7�P����v�����^��_�7�Ú{������!�x&(���R���`���<�5-�[��?���ʼ,]� �r�V�	���R�ՙ���U��Z�F8S�����ӕ��j�F���lP��xH�%��u��@�	uˢ���ѣ ��^H����b��r� ;<7l�$ބ����(l��P���?^�%B�g��T!/��W>�y���*&�1�5���q��׌P�@aP8���d�qq��^c�$� =L�z��Ay��a.x�ӫ�T�*��tfs����#�
��Ӓy�]��V$�,�m�����G��2�6�ri�h"(�e����m��?��@��%G��ಀ��b��������X��/W� ���[oi�#�t@��\�9< f�ǖ� @#�`%/�AQ�@���z�0nR���K��#Ά\�O�5p�ϑ�"ҏ�O5t���&�]��q������f�a:��x���N�6��T?�=n���4�iʌ�8��sU0���q�{����}�����)ِђ��3���%K"L	�K�1��ߏ�1�����|2��T��_�m!\��`ԭR�d�6��H����O���ѺXJ3��]ċ��Tֱ�(�7ʣɋ�6��7A9�	�a�2s���&��*ܮ8Ɲ*���T1���v#��[��jn���r�:�]��Y7ԉ�Z��$f���W�+���<�\_�D-l���W�$��0V��_X�'!�l�{��{74Z���O��7:a� ��{/[�\��*e���8N��Y�/��c�s��ͧ�}�=Oe��r�ʝ�%�'eP���O,�N�ax�-H�� �QJa�a�[����BIEInlswv�'�hT_�R�5�r��0MT����V���ӄX����O�Y����7�� �..��^����N�}@<�H;�R[��`��>��-�J����K9_���!�J�Z�Ս����:4��حY�a�]�HݘE�<�<�����7�G;@P��	р��?�#?D箉#:�8{�;�M.�#��Ɉ�hC2��|U+�_~z�7��6�̓�̓�Vr� û6�
Zp�֊�7uN�H`�zIehɵY4Z�{X�����?�/=�!wM����ą�c0�H8�¸#F�V��VM��2H��@Н�����ί��e�
�̌rQi����J�|A;V�WG�Iv>H����L�����r�<l��LRo���s�Uw똻�8j	�X@<o0oOG���Y�4a�ý�*����j�F�	l҈ �~�����I$��.:����x�#&6�Q6��8R�n#�c��~ϩ>�#՟M)Ri�,QU�d���;X��l�MA��D�!L:���O'��O)<dMxl&_X��L�:��j.�w�Jp��;*�ǥ�+`#r��kK���������SgՖ3�LN��N���>�@��yН9w9�kPGF�ȡ�q҅��O�p��z�/ˮ��y����-�l�?�A��M �����f�vz��DbI���]I�����ѽETNOÂR���7�J��
/'�xyĻ��ӠF�r��������&~m�����@]�Ѵ����&�\<so<�����:)kr]fV�h���r�C��lE�0�O+�%�(�X�'��}�Q�e�S���R�t�?��y�wJ��Yr��4��2뒔�ġV��� �1	���/$�-���G3��xZL3n�h}�&rK "��k*�r�!��ڵ�%���"+��Ow,�we�q
��jP3�p��xt��i6F�I�n�J?���I��<����e�5�tc\�-?XN��4{H�ʸk���x���lT�(/��{䒽�@�YUV����g'H���|A��R�f_D�(䞯~a�#g�}�ZJ^�P��N
��s𖛚H�p�Yx%��0C��t�_xk�7y��RF'�{\vj{;���R�O�9~kb^yv��E9ZUSx`*g�7A+��4F�|�n�b��Z�Ɇf���~s�JynS��Otj�.A�P�4��㛳�wۊ@�fS����##�xO�!4R�'����Xfح�a?�R\��8��)�����x��ր_1��6��'��%�))[;(T���s���q���?�#�Γ�;�U�o�'k�%���������I����Q#3��`;��kzA+O���t��J��o�^l�,靈f��H�
�XF$�d#�C��k-�Z��o��Z��0��%�$�F�\v,p�^�=����?Q�emMRw����K��XG���J��J�ᦒ����&OO�HR ��!q�Xc�����F}�M�G�*��oX��na`$<�o>�i��%����Jh�<��Cȣ����5��ؙ�"/@y�Y������jt5��뫼sx̍
�t�J��'	���Tͻ�\��.��Iz<������:AB��p�&K�nXٺ�뉎�|c���*\�Y�B��w�O?F�x��bܔ����uI��%A\8����Cl���X�S���H�'mˤ�#���reM伌Y�L-х�6�1:o�c� 0@�j�b&q&��(B@�٪��SH'�C��u�U$%q�����p|�����8�@�a}y����Jy�-���M�y�pb���1"9�o94�����6[k
x���2�-[L-<�� �^{Ӟ�����8.�n�C��m���S��2�(p���Ra��+�lZ�J� ���	�ג?����D��K�Q��k��[9��~N����7W5
v��b�$�ܠ��'��^b}�[�GC��D�L\B*7?��^�U(��؋$��m�zK�w.��{~�fD�!���r�C8]i3xS<�*�Ag������XA?���R�TNa�Q������b�<���80���fBgܬ�7p±�;�T'�ʮ�É?,y�{�Q#5�| ���-n��Q�d�#�v�ԫ�<�(4��\HY�^U����DY*����EN�&�rk�Cy#�Z��Q�	�\mA����3)����r��Ê�yi|;��&��"��O0`�wG�`iհp�X��b1d��<��C����p��ą�����*���ʙ"��C�rUi9O�c�z��!��^P匫�s�PLIg}�}�~��oi|�+'4p��u�P� ��)*�u�A�����t�[�,������Z�N�c8eщ�&PHI�Tz��x��2Fߗ����5�9������X"�槩W���}��T�a���*��:`tM���$Y3���!:8j4T�iN}���p@���^=B�d�O]���(
ܓ˥������I0���e}���D���S�"����')��m"N	\��aJ˛kK^����c�����6�(��Y����#t ���I���#B6v�>���o �S�}P����7�%Y1)���� M�w�=���GpS����Y��ڢ����NI��O�o�Y�}_����64�)8\��\j:&Z�b�7V�]F-�>�H4�Ua���bT
�	H�{�h00_��Ȩ�5Y�-���@�x�s�y~��@<������O�ݯm�=��4A<��=~s��·Z�4m�ݗ�������]^3N<c��ǳ���}5+n�w��5���-L,U��Ƙh�˷5�\@�y�p�L�fLi��"����8�?~І��B�I�����5Y�Ҷe�}����Md=n���m�ώͩ��<dI���f	�2�V�Ө�P̶����_��R,��!���C�����G�����̸/B���Ψ=Q��M���#[1Գ
gX���j��A��F~��.��ͦ�0!7�7f�ߔ�����83���D�L,2���� i)���Zb=�����q6�cRPL{ch��[lXeC�B���U<�G�Pp���ܹX���j�c�kX��q7��1�2#���i��f���a�(�^��F��m����S�9��㞳��jTD'o�D�b�ю�5���j�]���H�c��+W�I��vݛ
3��~	s�hq�h�4 Pr�QZ���*h8����姵a����Uל�ɱ�X˨ c�o�<�*癅����O�9����z���{�d3�އ#�w�Ь �>��@��Ͱ�
�ˆ|}�|�ٺ���=7r�@���`���go�LR��};�4�n$�#���$�ljF1`�[�I�.c_ݴ���ϭ_�v{����'�
+I��?�6� �/݃e�*,��|��׋?�z����-,M��tlX���~K!lC��P���f�8��m��=�
]�):G�J���\��g�\~J�:M$��n���z#�U��*�cF�q��Mp0,b�b~s�tlGr9
�%���3�D���t�~L�����~�8lO�-��F��k�(�����)'g1�3$��xb��d�"H��g{"2�$- ����C7UQ�-wI�ɐ<�>`��xG����׷��j����� �J��;�m:�aw��mx�B�c?��;��6BUj�l:@�ŷ�%U6���&5����Ǹb���^���]*��߬x��U���<8�t�&�.Q���\Y4��o��ܞd)��)�L*�����Hk~
����dM�H��S��+�7�,81��<����gZw#AG�m�~� �7@>���"��{~���,�`�u�Y}������%�T�i��r�e�(��|�E��`��g��.8�THK~�7�h�˹揦��`Z�g�߻�&^-׽�e�.�5��o�8�̅ﹴy���ȧtk�2�8ΐ��?:�>���E�;���K�5�Z�4l|G7`��:Ն7����`�Ɖ'�#����Ţ}BE�)ee�z� ��t$C(�о�X6E�%�=��dCh�sk|_n���I$^W����j¸*�՟i>� �����A�S_�=O�tƧ��,���O���̻����:��G}"��Z�'�i��!�=͈򪏎]9�lm�&��Q����.OQ��N2�v��I��+�}]�<k���i�%�J �1�5)
4�kRU,m7�A�x�{H�,`�	��W�?�=�zу��@��^�?�|�-UP=_��_ˀ��/�VĹ��L��Y�����'�L)�8|���#�ߟo����b����-K
�w��"�������U��G�����'���(��<��	y��,��Wfu�w�5��%1?\�ؿo@u�Qc(X���L�$)C3�X��2�~�N�(�y���r3����5lf�&O�X$%��CL���J�W��5i�(�=b�,�㸿S�ߊ�$��9�#!qNjV���*ws�F���_�V%�Ǉ`���`M�q��E��:��h�ӄ����r<\2� }%r���4��aB��e�7��ԡ��(�P._K+t~���m�/)�*�-��td���q*F�O��su�� �����	K4'�I����pCY���KX1'Ӂ'�.%Ĭ)5��t�^=��|w>�Zx��4 �84�#.7�a�Km����jO�v�@ed�3Z�����
<�Zz	ׯ¼Z�Ig��a{�sktm,Rt(�Pv���T��*j�~K��; ��>��vmym��pƵ+Ԫ������<�p�
[�ʒ�Z�`	�xф>X��|�����:M���k=-uDw��)w��%���,��dB��˘�����t*K��؞<;��ߢ��E�t�=}m]�,����Ջ�7(�9?+��VT�Lr����Zi�I�3E���<�)���*$2^�WÅ�|�oؑ?lE6��fy�ӤcB����ŜZ�ZH��+��zVTN�2��f_f�3�dz�}7���8d��FNCzUg�����܁�W6���޽��E�ؕ(�>����b]a��kfT�� {�s��	���?�P��2r}C�͐{e��B��v$ln!�;gY�<����� S�J�x��l� O��+n��_A8�W���)�5�������0�B]�@#�h
ǖ��/u�N2�N��寲 �p?[�1�k��BG�Ff������KtT]�K�sǝȨ)�v�X�.dF;��BV�9+�

����O}h��ӏlW˵���\��-Hd��C�z�뚥k��G���T�0qw|�����X��������V9���1s������)ǳ봩�� �S��;�i�J�W�mAN��)�0�uL�����]q�k��U��6�93ࢾ@Zo�=u"� ���zj�D�o&H���v���*�Z�ܤ�ˀ�ag���!������	�[.>R�u$-|�;d��.�oa�١��Q��+��
�8��FO5���lb0���'��!��c��)�Mޠ
��@�E���^j�!���,��Yz*[:�1��ѬQ��}}[���v���(��
]�sE_[�ip~㪘Z�����Ԕ�qZ�����ˡ��S|��gutVփ�!c���lKC�|��P�)�+s��
���͕V{�}���Y�B�W�en���-�|d�bo�. ��_A|�i1�;�b�d���'hOʙ{LY��d\�ue"9x�T܅��!!w8y�X��lWI��0m\J��6OuL��`ޗ�LV��������B����ҫy=mT0�.&_��+��i|>R���b��k�5[�|��'|�>��([�E���)3,�.��� H�8S�?��rt���}F��6&xs������E�} nsl��V8PmP�)���͢'�E�A��W�}�j�*�$oJ��.T����l�Ď	1߰?Bk�����;�J�H}�Щj�������f�QzH$?Z2�M���s0;=Bb�����_�fDo���)=Y�.-�n� DA���vS��G�今�C�!Ȕ[���z4�qԾ& �C��S�7F���!G[j�0�����r���,nw�W�Y��pg-<T�3������ ��Lm
��!�[�kK��H��� ��);I;�/%�*�KU�"�
���6u�q�y�!+��׉݆er��΂�oLY�5E�K�)'������fBK'3[�����'wY�: ���2oM�,��a��y�SG)~��C���imK��9׊I���oZ���V�s"���Ǳ��nʡ��}�|��s����2���%��b_��ğy�M�87���hR�{X�X����[� �A�F0�IB`�2����� �^�rA���?�0��y��ݖ�W=+G�����4���m����X%����
��/n}&�l)E �޸���usJ����1�_s,�/p��L�՚K��w1��%�ǟ(��j���s���k���7�i���;���4��uŀB�E��m4h+I_u���'m�=��N�4V&W�����}7$-|�a�V��<��RţX�|�'�I�;C�5%Q*�g�o�p����< ]�H�)�@9��cǉ�|�&]�W	Q�2�����`{+��
�(��5.v
�w3r�����	�����}m�JG�9Д�̩�[1����Ǿ��i�Rg����wX�̡�I:2o^CTh!���<1��$	� �j�aM��2�`�EvQ/&m{�1qܪ~4�?�+�� ����}p.���z��n���Vه�Pd�fh&=�,�m͙��2��=" <�"Q7������dN������}8�c�C�&}Jb䤐楫�*�Ц�Ր����S�>��.
�.m�/~�ce��%ƚ�tk9�4sn��.��J/M�@��{]�$~*�GҦ`���
K[��A�9|X prSN�6|"<�k�F�G���v�k��gPT�y8��ڷe���MkP�
�>���6��Vx����:ڒ ��y�����Y���ŉp�¢R���F)����M����n�D���^ Z�]���������5|�?�:���G�n\k��xC�T�c�S*o��#9^)�w�7���P�x�􃪾^D�l��x��)s�sāgb�J�јE5��� y�,��Aei�,���LX> ��\�@��H �Ɩ�bo�Y�EtLAG�䳟SYPP�,<nTH3�O���j]RG�f����RW�S� �_YR9����Tu�=��2q�2�JLHK)��_9�w��Ts!E ���-�(���d>Z��7��pu�d��_'���-��l�Ң�O�Lxs�D��\��u7��Z�em��WP k��\WFR���k���[�|8�x��Pr�{�Pt�!��D�#�%E�F(��x�n�B���V ��s�:y[m�?ɼ؉�T�^�G���N��g^�#>z'�x?���6��~�H��.��%uh� .�7C�΋"�5V��x}����m��h[d=��z���X�hC��E��.�^$N��<{����͕�4+����M!�}p�ZZL��_��A ��CQ�f���*�0�9/�>:-J�u�E�����Av�����y��N�_�����="�֢(9�i���F7S��o��DS�T9������C�P�]��\4{a,�2�ͪ�U���t1�w�*�������+>�t轂��N����0<�RL����*��a�)��57�m[�bw �C����-5o��G��zγ*��|��<P�i���'��K�р�d�H���L�>[?��}a�y��/��܀�`#��J7���ߢ �%�hN���q���%u��#3wo�y��3�Y�t��ͯXm��Xi��;DH1��7�$��5++���D��%W���fM)-�/5xC+&)�۰#l(��$4��	��ۢkb�� D��N��G�'�7�zֿ ��I�k�w�>�lXEDX�uj$iHg�k�^���]Z��_h4	B��k�v&��S��8Co�s�!���0��*%/�� �D�����|����0G�hO��+$PЭN��}�7�����A�9c�Љ׺Sc�2[���6�QK��(`�y�w:,"}_찄o��/}���~�J3Q����^^c^�'lc���r2@q_�:x�L�ΓS֎����Q�Ö��I�����n8r��&�T��Bck��3�w0ٷ�!�B��Q(���jF5��l9�a�X���R�pD@(�z.��>�|������1*�WL���?oT�+�Aj��`B��Ϧy�2�9�=���L��ܐi��P�mQd ����)�����$�
>,�������À_��������Z�"�u�!s	���+�ᛉj��q���S��Cw�:���\��>e����	p�רX���Rbt���#7w�&��R��#�d��t�s���a
9g�?���A�Ol:�.Uѩb����I��X)�S�W!b�y����ח�F��	@d0x���/�A��]Y�Q�JГV���$�-�cz�j��6�#�K�3j<�u+ũF�U�SEV,,F5�T���Wիm
÷ T��(*vմ,�#������W�^D��E�ՓՋ���hǪ�=z�b�@F�B�)LDW�=&]X#�C�c!w04����W��Q�c�T��5�kQ)�3�d�}�g��0X��)�A˿�����������e%�)V�9��^�w@��W	yԷ��Z)��"�%��]n����r7$Yst� �����qsՏ�<�xTS�**�4��GV)��X��Cq舯|,�\`��X
��-�f�����Rc>z�B�p`0�wlw��_Cc��"V?4� 0H{v��a�T���cL�_oj9�o�!0i���ӿSkq@{��0��%%���\���}�2��zPF�
s��6��1�tU��xi�3h�tQ7�L�����jm����4��-�՝�����Qa�
�mfw)�\f�b��	�j ��9Z*�UjV++�@ހ�[ѝv ��t����۝rf�Q�"�n���{UQ�liyT������]�*tL0p�����@&(�\�'�:ŀz���34�,>+��!��!P�>{R��@l��1�m����:�9(�=��Y��ӚƔ���g�
+��6��TT_��=p{�*�d�Y�J�Fy�l!Br�' @ ��� 5����ʮ�ZT��U�U/nV�,W�d�x����k��j��-��������@1�
>�E�S�[s?[/M�n&�e @?7��~9����X��^�� (T�S���0�r��c��*>���T-��=������xOFX�D���%[��}U��%���$�ܕb�e�J�\p�lĹ�V��/�W��\~@�"���?�Xj3s��ncc���?f<����&]�}�mk>]xI7�o+uU�~�>���}o˺f�L,F_i��7�5T�ÿ���04��r������Z�Q�̴A�v�[�x"T@k����ًM�v�f�YԠ�F�PDIDxKɓ�(I�6�J�$0)�v�1�)<����1��EE��5����(�,�)�(�q��`z��R�0E�N��l����.��P�^���=u_s��Vt�.������$�AC�~Q�vl��/���ըݝG~`o�������=�E2L��>ۇ��+������Y�<�~#f]��lI��v���/`3���|M��c�ȅ�~`�lc -8�zOTN�O�Q��b|��Vo�U��t�j�I���_r.`h�1�gt���h�ͥ�CK�EfC�4�]V����%������Pg8��R�݁y:Z�f�Egl�9���{�p.�L���aY̠��"�򿋼��j}�3x�	,H��1et�d����YpN���D
��\ߙ\$�W�A�BuRFM��5��s��?ݑ���y׮�$���E�`� 󂄿zr���6��nF�S���� �~2'I2-8��܌C��m�%]�������1P�>���B�(uQ�߸�Ci�0'��%=r$:f �W�{�^�x�Z��A���0^���
F�zd ��x����8�7+A̯;!tՃ���4@��7cy&��L�� �A���"K��A 3��H (�gHc����c���iqh2"E
�.�?k�oP�6n�Bpޠ2�&08��Fueu�=����6�B���o0�dgا�U�s��Ib͚��亂�e,8|=���-P�,�:���h����Rs��vxڄ��'^�=,;�p���\���B��a���A����id�"8=M��b�ԉm���b�I�٧׃0�E�Dl����%��`.�lh���P��3Y�T�t���q&�(A���ֱs�@zM.Q��@#��u�V:�m�ó�E|UB�w��!�F�/5ءF!$е��5Gp������մ�b
Q������=P0NhS�ȋ�X��U;ZR4K蜒��t){0�>��/�0�*�[�R|�������L Z��JU��Ęr��O>L/��M�"�Ui����k}~U��'o�P{gq-T�6��1-�n�F�B0�&��s�r�L�M��z�qG�$����g�I7ozL��y�d����4�v{����?��^8�O�S�~��|�P5�]���5J��s���n��#l�鲓W`���{�S���uՃ�:|��|�!u��"�+N}���q
攃q�A�tt��#�w4Av:w,��G��Q C���cέq�S���ʲ�D ��3'��RmU:߱�ItS?�t�ӆ�(z3;^�#9�E��;^'	�G}�զ/NQ���|s�y�<'5R�vHv�h��2��m�3�ʟ;�;g�lCJ�1���ٿ�g|9̣�����۰���{����AN���no�R�����L���qh��kі��/�k�vP9D,9��n��ػ�Z��~~��L��e���s��Z���������P��鼼	�BO���E̪s0���EЖ�XG��i��ܱ�Gm�\+U�l;����� O˅�n+�~��/3����&0��>���IQRn�@������;;yiA8��ݰ4Q_x���6�,Ӷs���`~gwy{��%��S�QJB
�by*l}{4,�X�T�!�L
�.)��]��ͺ|�]���~"���_����a��8�3ƒ�p#�A� 8b�����W���<A�9��/ds4�*H�.$���1�.*L��EPڍg��)�q-z�WJ���s��5��2�'V��)��th�t��uW�b",�o�� d�`�~�C�7ol�P��i/N�7���@�%1�Qy����'	�����to�n������O�SX%�x�����0yH�N���� �`�r����ؔ.�2ـЭ�p<N�r�*g�G5�+f+<�Xy�8�������n�*d:Y��(�9.��Bݩ$�g��3i��{|FQ+]_Z�ݎ@+N��+�a��϶c]_�q�b�i��~�W!8�D[�R�0�!�#�Ag�����L��4�Ռ��a���*���.	��4�o��$��g���=i �)tT�.�ǯøk���a��D�� \�~ŃQ�%�"@��a2*V	��\E��o���^Wp(�YDS��݉z����}����/9����T�(k��2z)��W�8� [��F�Y[�	Ⱦ������QH��_|��oy�y	�����O���a�G���������{��{(+Dc,�wm h1)����ri5�<��	�I����(X�H`�Tls�\&ē��Ņ/�XU��2M����-����/	��Ωu�/�uhQ��oo��$��YǙK�ɼ�����9(��$���8%����5��Ts�)�5n&����>+�R��T7�p�_������>�b�Vk+�����&�'|�a��%���$N�l~B��@� 4�ߔxZN���P��� x���އ��qʜcN�K�i� Q�vI8DP@�cO韁V�D�o�M9I���٣Y���,����0��̹�
�I6S8��ץ�8���Խ����#���Β�DS�wx�P�	�2~q����T��Zʹ6�
P��&n)����8��M�~����ȇirzp �h��zO�M�z�8�m��W6e�����@� ذ��
����WH��^YE���+u8q�M	!D��<jMp,�O��m�"Ң����-t�n<v3��Hи�v�R�_���e4�Y; 4RK+��(�"�r�/ǁX�\΄$�E�}�q6l���t9)%d�"֝�V���io�7��/�y�>p����4����u��>Lm"I�>y���)�逼VG<�3�Zm��un�Tm|�C��?ҽ �n�]~$���R,��I�����2<�6�E��a]Z�B����M-� q�z9 d!�`�����!���4Y�%�x"�{�͞���W�</Ey�?h��j���16(8?q��VJ(��0̒�6����o0�GK��&s��d)���e�l��Iѡݰ�LÓ�ҏ��mv��`�G+�g�QQhcYhP<AǪ"%"�ˁU�����bB2e�5m ZV<�vY�Y��S��L�_z~�n�_|��i9jVE��*��^�?M�ĉ���F�n?�����\nV��"0lӔ�Bb]�u	U��\�p�c�d4IE�Ӄ��Bd+=�.#�	�o{]��+3V�lHu�_`��1�)
)���s�nb|��h~�e��h���9f�e����з\B7�G �!��)��`��U�J��K�i��K2s|Hl���1�q����)��U��Q��UI���!ʢ�<��HGDY��R�Zցk�y�z�&��֚FG��{�ݪ���L?_T���{+/�/IB!>�� �*���|����ܐ�f�kP�e#[�Lh����z�$���O
	 rV�s[n� D��vmt:�+�;r`�$�We��Ǜu�aQk|#C
F��9��L���ll}�I�%蚶���i9/���q�o�*��뺙:
��a�F÷�5\��r�����_��T��e]dCW���s���ʘ�霉'�&�!�l��vY��x�E��'���#j�Z��>�=Gy��3ko2�A�S���}~���ܭg��,��5��%7�sF �^���w
���5,f�^S�;�ȣ�*5
��ٴ�H�;������V|���V�a)��q� 
��a,�q&<rR�L��߂J���m^{�,�#�\��Gt	Ew�����#6�}RU)��k�1u��X*:�@��W�w�,hY]Cc~�9�i4̓��_��vr���b"��h�ϋf��Fo�}�)~����t�1;&��ς�@o�x�hz���⫉:g���@��hPz�ࠬ���K��|�\����k���6�3�ŧ���T�m+S��ȶ���{�i űP'=�uM����5w@�������6���vD�<B����w��x�$�8b���ՙ�I[��R��*�w��ӄ��/{�|qt�A�ǉ�}d��:�U`#��S��`�}������y�	��`��؝Gr[2eL�����Q'<��C8�o�:�xq(�.�~e*�
���M������:5�lN��\��o?�<��'^�6��5�����1�Ղ��m�o;�ǿ�L�I��H!JʖmRGؙā�j�r��fe�mY�qT��$����)�u�����"(R�����8S���(�H?�<���E8��)��ާ��%��tO7����F�L.�
@=}�� �iiՔ��7�M����#�+�\:�0j��+).$�+\���=8h��j��r� �x�\�c�ϝ��Y}N�cS
�-�4��mr*��e��7g��}3Ѵn��r���7�ˉ4�#sK��J�[��2?l1����%gc6��~!����t#!L��,�������!���c����p��3S�2����q���_Y_�[+�o�#�M(��.D�,t��ЩO�U3#���w��
�a�)T�����(�h�SEQ�����֕�ϱ�%V�A��B�>���ӿٗ0}�V��܋���6Q�~CF���$�����6��1������jŌ����[[��nc�s.we�lz��C��$d�q����K��xT`ݱ]���ꀴ�Đ	����2����G G��[t����ڜ��U�27��C����w��ō�8k��U,�R0�/���<[ς��b����Y��Q&����M	K5����G^>\8��NAv6j�.�{YXO��LS��v�6eP�
�f�t ���sDl��٤��9HF�!�e�ՔS�j��F�U�0��n^���0$��m/jUh�0:y�w�e8�Săg��Ѷ�k/F;h{@(s�
�<�Yؠ���͢��V��-��������r:��i{�� {�2-�	ۿ�q��8Bt��оP-��U@藺���o������y:����Ԑz���L��D�����]��"���כ���m1t &ǰ J�����4�r���͝@��%l�����z�-���Iɡ���\|�D
^Sǵ	��k�Uf&�U�K�t>����z�=��:^�Ζ�G��v�؆Nw�K�ے]���՛>��r�#d��g� �aW?��U�-�����|��-��d�D8K�ݾ���<Q�|�Fž8���vm�V4������GQ�&�J�Ut��*h7h��Iۻx����S�����ZLK4k�'���}�6��e�2��<�jn��gl<o���GX�S�q���C�`�������s�pU���m�:�E�|'�L���8%��� �`���{j!�֫�����ac�;���`�E\����~�Ixg��5.%%_���L@^�w"jܩ/{Ld?�Y��@<�9S����b�m�ťo�?1:��wU�pdSR�3 �C`�^}:M`����O6�o�{U��iI4Ų2o��޿-Nu�ɳ��(�M��-*4-���L��<Dg~�΋���%��@��$�#U�Zb�!�5�h�d����:l�'&<A�Sr�B�QK�dG�	ٯy�R�,�+����]�X|�j�ߣ� ���02�7#}�z}�h�Er���H�88��i)��IZ@�~��0pW륩�o#LS��\�.	~�FD9'���O����!�,��Z������^UWy@�I�D����c4<幤e]�]��@����F�D������bo��@w�M/c@����Z�=�%uM33��v��%7���� \�c��a]i�	��@��7�)!	�)��ۗ����\���59WO���4R,��A�I[�t7\@E�@��~�����}$9�6��M��B������Hk����.���j�f��I�{�z�-�n��z�m����V���~� ��0�ҊE��թ�x�bQ}�QJ���4w�{�o
|��x
)�+�׳,a�@�@	�-T@%����*��K$�Ŝ'*5��|���O[������g��{�9i�6�aT`ʙ�G��G9��Z���-{�*���!5vq�%��ʐ�41&�ᇜ'����2B�?z�/eP釅#�KFE��)��ӢN��&�6�;��3E2�r�R:��D�t	|_�sB�S�������u˶���B�ִ�ҏ���Wޱ/��Gs6� C��\\d�u�~�C�y�5�_F��Lż�X������W�)7��h	���^W�!�r�D4J�����fe���E�����mI>�u�Un��-������s/���E[�W�I�#��P|Tm����نT�H�3��+0ȟb(�'5�(Q�wP'/�R,8���Cb�
^��҃O,7�u!�ˋǸ�4��[Y���D	--�I�%���� '��'��$����3p�]��cRKl���/�|!F���D�o(i�>_m�j]dV�:v�b�|S�1��{�6n�{��	|XG"�3SpcC�V�Ɗ��JKLdS���U����,�ю� ��*y�]�L�>_ޫZ��I�����iꦰF^@�e��z
֞?�v�R)��\޹�����7_I1���k�C�;n��W��tM>v�@
��u��#��2���%�ȥf�;�g����dt]
�3���eF0-	N�ρ]�UP�^���5^A�j�	���Ζyz��9��4�-�-ِ�����-B��:��<`�s rڔX�|��s���ww=݂K�ij�xQ�+�τ��������*��o"��|tB0�L7�X��אr��H^�SR]ы���:/��~:��݈�ݮ�dpδ�1�z�0rc X�9��@�8�1�s4��g��JO��^d4��ĨA�!���{j�S$$֙�ꌨ�Q�,�8���s��T�S0��iM��po�Zb��I�e��=��U�!!��*}��["�5�.X-*c�a*��@ؤ�o���%���j��>��؜�y��rPpt�yb/�8م���'3����� 8��r�s$����2����8�ޚ3��Gw
/ѽ�V�0�<6�9x%-��(�eg��Pj�r�5
��ΰ��
��y���'F��.Z����`�)�S��c|��mtu�[�.n;���3�\�|���Jy� u���5<�f���zZ��Ab�o��;��Y'���Yv��툾Q\�����=v�����OHЬeBt�\R<�Ơ�O�;c�U�`�L�(��&*M}�$o�>�8j�'����zH���h�5�}��d���8A�ٖ |!G�/c��L^24�ćT��kΒ���%wv�K�pgB���8��K��@@�5?�r=�1�c���@wr�}�?�l�߾��#>-��A�m�����;��"b��Z���vr)�_�x��Rއ��W���"�;�`Q^��ŭ��+Sq_��59v#T�����<�S�5���k�:��ig.ݮ�x�B5���ڗ��#�����~�"��#� �S���B*ˌ��§�`]�3�נbW�ZM�L���{�E��Y�	����u�hJ�$����<�a@o0U2�Ҕq�~�Cs�D[��E*�I"��7�U~����ik@�iQ�A}Qԑ�&�1Ϭ%R���U��-��u��y���E#h���W�����Rϐ :9S�U�4OU�G�""6�|���%������R�}z�ŸJ��4 �nx��TF��G��ɉc2� �d��S>�4X�Q	_��!:�yD|f��|~�+�[A�\���7�����8!����l��C��Y��)\dM�]�NOD*�����
��mUʇw_�,dӈ~��Q���Y�v	{�G)�"~�$��nk�"fM���@����.�V�rm��D��{D��p�s��c��
��&C)�s�3�[�-{(ə�*dz�>�4n��c�T�:?�v�b�qO;��E��j<tW�6;��\�G?�]C���jA+s������,`�TlA��/�1������!���5��JF�r�J��9K5��t!MƑi���%���ˋ�@�d\y}�b��vS�I0��S����*D���s7K�����J5��Q2�s_���B��xr�@����f�} #��Ki;��$t�)�@��W5�8~�b65��
Z��̴�6*����E1�$F�!>`)�EШ�,�961
���H�n*�lg>��9��`jz:�H6�\���7��kT�,��稽�&v���g>�V/�j,�m�z� 	sO,�>$�f�d��7�s��u
 �J�^S�X# �60��R|�x�@�����2����[�'�R�M����ROb���FoW�,m��O��ybu�����J��oo�C�cl9^]��\��|�}R��Z��b�X57�g�<��x��+���/����S3�K�;^f}�ٙ^���ҧ��P�2?�O�x��;�-�RJs����DH�'������k?3���=�y�}]�s'1�K��1a�K�>��a�4`�&4�!_�\��(58��5>���ܖI=jS�g����M8�2�tTbbʔ)U�e|,n`�P߁f�Ӈ�&�4�!��1���BկQ�<8�1��&F�d����ה�D��,�9+Es��I/��^��or�e�䠺;�<�uT=�>�0�������?���z�Y�1��oA�so�M7@ų�{!���h�������9T��3�!\(�Q?nv�hV(�R�\��=� b�����M��:�GF�D[�\�nK@:H�:D#u
�� |Q��t�E
w��5���d��FԶ�m �b�,Z��ǃq@��q�J�b�;�Iepx�w�P�~����9c��ý7G#G��I+0�p��D[:l(=�����b���z���N4w�}IW(>7N#�Bz����}^'nE�C-��t�L�����u-,�6u���&:�W$|��>�S��خ�e�{X��aeVّͬ�>cZB`����%׺��h4�D�����6����f��M�+in�:I�(�mCilhb={�V��#�hȠ��vRS!�1Z)ʟ�C+�8��b�[n�5]~��CN��4�Ǖ���ۤp�t��y:����8��`��{���䗚�5������	��|�g	����G�v��Ala>5j]�	
��y-b�� �ӡ����O�L�Wq2���q���w=>���%29�ȧ�}�)o%Lr�ރ_���fi��rݜ7�\!g�5�|iP	��$6���d��!�y�haH����H�֮O	9ϒ͵~��}�մ�
���nEG�ho	^i��[��'d�O�K�T�sQn��D�A�7��|�)���ċ�Y@�`6�v��#�V��s@eN�"�3�vC��hi?"X:~ݖ_��<p֥���\$��}��?�e�e	�V�1�PB�٣!�$/�%�[
|?��������I��5H��$��w��;��~�0~���{O�����l����]�<�dZè�9��l�6k{�Ҝ��[b����2;-�a�mTD�R§���o�4R��橕���Wm�\W��9TU d�� �U��w��7e�;�"�Y=�8�f��~�Aٶ�~�v����]ג��.'1uAq�������-� k�f5���;)D� ����(��C��iO+P��F�Q��J�8�p9��찗*(V`�݄�+��vp|��Z�T��hwv9�=S/O�ų{+1�B�����Z��A0ޙ�T9�z�t���n�h�8%�cu�rh*�٬�U��8}�f0z�!#>`t�`�����YQ�3O��0��kO-��G8!h@�S$_�*��O[�����3h>^.ݛ����9����h0$��[ķ5,כ�_�+����w~�eF�:F��F����U��L���zf�v!e���"�c�Q6%��S0Y���C�x��*�_��},�aR"��lF����7ꜯ�������� a��BV���=���G"�[1#)�O���79��}�~jw&08�VX`@q��E�,M� ����!�R��EU��;r~ :k�9���=5�[��M֋����kj�k$�Ԃ�7��� ���{���f�i��x�0�� �.��BV�߿�>�_%O��`i׷*���q�3�E�2���~���K����C�9r3sѫ������5�Z�VH��Nmx�X?c��qǪiu2�c�q�l��?�9�v�@�t�W����[�Y>E�#����@��� ����q_<�����A	�q�͍ǮT�4�Y�zc+�>|!@��;�354@!^q[�LO�EmCf~�$��t o��Ӯ���8��	
��`�A�F2�� �Z%�%�"\?9��E��!Pb�7��I�m�L�+/�U89M�c5�����He��9�F��[Vh��X b�_77`�Wh��$���R��)�A�=	ǮJ�����J[�kO D�b�,'?�@�Z�I0鞧$��Jt���H ��i��{�)��᧌���Z�8Hm�-���X�7Rb�C��5�i}E����En�EXㅶա�\')>vi��శ������Q�k�$?r��!�MpyxRZҠ[�^��BOʌ��06��]ǒ�H�<X��5��6��&�t���"�n�6%&N�@�J�o��=�u)z2B�S���~l7�Cgo$ e�RY�vtD����T4�.5_1����46�~?�����ʒ���J�3)��8.�A��JD�m_iq�1�v��p8���fY�T�e]gn�ux�ń�n������*��A�DGBg��w-�w���tz�S��`Nt�+6)������;�N�=?�a��t?	Tv.@8�6�ag|�>{6/Fl��}{���oN�<W�l1�>�Y��H"� �bA�1oS �LϨ��yq�E:.�-�ǳ�4�i���$�������W�I�xO��f)������MY��Ӝ�|��������}�j,�`0�=��*7%p�q��V QΦ3~��8�>}�㳚�n1H��(���If�n��u�,���I�L�!^k�bo���kM8�O����7�IH��T]�K�D��)h<������0�j¨ s.](�	1kn��Ƥh.�y�c!�L�	�_�^�h��[�݁�a,�P�G7?�y\���#Y�+�h� �i���~B|I����t�:U��3y����ZE꠳>^�9��֢��>�Ïl�����a���V���W(��c8��j���ZP��*s�a�~�T�o/��3VRx�I��ˌ��QOY��d�B�@`#�2��~�ecןۘ�TJz� A厹�PByLu�|ۦz�e�������^�G��{��r$���/��/�]�Mb�f6:�\�}�s�3�y���4CWPJ��O���(.H`��˝jbT7Y�������� ��ߜ����<R<��	L	��lQ�����jaO<��\����G �=1�ץ�Q\��ݳ�c4����q�d�� B6@�W+Y��JG�u}Hq	><��P�Yq�2�`���v'�V"o`*+��-X��,j��,�\�����N�E�mn �7Tk���#f���NkVB쮡��T9'��&.v�-�9S_�*�!�`��]%e�nnԝXP8�iA��2E�:^g��!7ƪpHn+�)1����C�w�cp�<�I�*���A��
���<ʴȕ4�6��_>�E����]Wp��b���=�.Y@#�'5I��^el��^����_f���*�M�a*x��-u����[t�c�u�y���ӉL���1�d�d�u��f)��+�7�v�<� N��O��9�%�N詄�>u'�.���
d�mg� ��N�2��;�B�w(���=��.u9��	hX��n�+f�HU8E��6��j�]���9 �4�F��d����FT��Z���%��+��%;����׼Z��I!����/���۩j�<j���a[(�Ï{�j���Ԍ�b@rξ�^�-)4ׂ0�������|���_�j�d��]Mh-����V�ӂ�G��8Հ�:�J���/7B��Kƨ�yQr�r���h�'TS���xr>n;���P�"L0l9�
t�\p��ZB�qO�aʗ�|�t��F[?�)-4u��
�S��z~���{��+��%F<���5l��,�:�W���3��'�A̸+,��M�v/�Νh6]��AM��xY3��_p74���V�ɀ����1�@1�w=yD���jho����c�f[aP�����.9�!�g�N7<��S�O�c9FZ�C�M�Q9�������肪��� �Mѵ����$ �S�>A� �J�QO�F�1k�5�����D������)w0@z"�wb0�&N!���Y���n���ĭ�$�7N܍�>��S@j}�`W�F�bZ�����]5�Tq
m�������}��'�+���yY��<���ʦ��!�Pq�$�d��m1��)%�&~0�ےw�"R}F�2�k�C?l�	7>֨������*�V��1�%p�1�9${�(RMO͔L`�W��x��ַ��8fê���@�,3Kj6[�_�<��*6�
�u|�en�i\�r.s����j-��8��NDz=�'�0J� �֊Ah���"*Pu�- �ú� ~l�qɣ��K��k��E�_����/�ά[,�V~6��f嵶��+�/v�GJ���k���4��6%{I�&��N����췹�N��|�׍��aF���B8��\A!�|�X�'h_�_%�:!'+g������*K�r����}�g�hQ�4X���f <A���װ�i�Ny�D��^M`e����'�w�U�{0�"}�T4���+~�G�3��O���������#�BH������Sf��C�W��ӛh5CFG_n� �綏p�V����$��1�r��H��<=��N���>ݪ��x}�~Y���ZS_>�in�� 	��>�����g������nJ�˾���A�{�����<�a��i��/���܌�,K'�`�!�z�*�YI4g^��(��\��;��/�g�`�98���i�j�����cF�H2#�m�N�e�7m]�gi.�ad^:c0�/�����=Od���\�S�V�����S�x�G��Op�6�WE�����[0G��9v�oZvs)�`3$А7�<�	8���D���̎��@~��C�*���"[��a.���!D��T����*���Goz�Ԩcׂ�>����
�����~�Zsv�2�,�rB	d@_�=u����9��UH079b�WW�)r_*�b(�V>��KwO`�Zeb����uf�]���N�F��z�˘!������k`[q.���FO��8@!��H���	�ϐ����m{1�f����;9~��£��9�q
���%C\6K�r,��M�F� �ِ��Ћ���b�1P$��e�}nC�I:#��"��[Ê_��䊒]5�@�\ƃ���"����L�Et[k�����>��4�p�i�~E�"{dy`׬����ˈMx|�6�kWtV+@�9�z�e<0��������õ��M>��7���yi�����7c�x��<+VM��d��,7�I0tOH��)E�(I� �p��>�&L�x��U��6� ������=���?^��������Je��]��lX,��#w���x_Rv���I��,�y3��<#�w� 
�k�/�:L���p������?��|ܫ�>�}e*?��,��8ί�3�b�k�ٮx��"�_F=|����al�f5)�K��S6�b��Z���| BJ!þ�9j[~�_�ʝ�(�Nx",�m��&]�!α�����ҡ�Y4�Q�x�Sa�n�%��<���lK����J���̧B`��g�0dr0��K}�8NA�g��~�^�Ǚ���Mxk���Փ����X�fh[c���7==��]L�a��I���*��tވ72%Ԏ���Dn�F+��\��9x"�R�S��F�U4.p蚪x]4*�`��8V\^gN�W<4�P�K=q�J0�H�;�'RY�BB	���0��E�t����t=~Kҧ	dU\�A5��-J�lnE?���S��ޔ⻑H��[�Q�(��br-�ނ$��\޸QiK:y;Y��z����倖���셋��q�kL�)�)6��>��D��[�o%Rm\T�y�sG�}?H�R.�X�~�N>x�����E��z���Ht�p<���}^J?"'�5X��-��ǒ܇f�|ھ�4�Hg�����,�Z|�;`h4SY
��xi��ct6!�!.��'�J�<9Ä`�'c�!W�螈i��Zm)x��v�H@�.?# ƴjÜ�=ߢ|��t0V�f�țj��X���?����q3s�>���T���A&�%�X:_�O�J揈-� �/iH�T������5Z���[*��F!t�-���Wm5R�і5��7�Z����_���|b� O��8�3}`��k.�Ij�!l���֩ȉ ��4T��9n�
��i\�v!���,�)0}�A����̴��ꤐ�㱡�R��V�5��� Z������Ț�u�w=��^�:%^j�W0���0/9��p��h�>�kAy�5I(̸�v�t�E@�_����k��Jļg$�c;�¯.� \ʧ4]
��9\a-�{�a��cʾI�j's�e �
zp�L�*o;�i+�-u�V��=hd%�|Y�i��FS�2U���b��`z�$�b�bՏ��넔��w�(�q���m�����"H��$u���<@�
�|_Tk(�Z�����s�vD�C����	.�|y;{f�"��)��ޱ�����N�q�*�@"�>���[l������Ѱx���m1m�=��1ۯ����ˎ����H��|����Fҕ�O�A��{���z��}2����L>����t�#B+�}���K�m��Cr\��JTú�~�èOn��}�56*�2!R�T'��x�yK�Wcp��0�53����\���cn(��΄��?�7u�;s�"`�6���nD��2�)G%��P������̼�p����.����]{�;L���U�|�f�Ly*7��M�>M�6�~��1_� 8�͓m�QcǭFI4 s���ؖו�n]N�}��Lô��AȚ�;�)�'�j�����,��8b>`�Ex`u"��آPk�Y������ێ&&�̘o�?�u�����`v��AӎF�F(C�����9S_鹜ǩ� ��Y9���g����2�,��K���0뉞$BQ#7Cc��yBf	�j��>/%X��=�g�Q�H
�E:�!��>�9ܥ�'� G��5:�#HCe��hn㮵l>� �?��������V/�tpէ8�e��u�C!�q������?g$��IKpf��t�J���S���k���cEt���È�R���j���<?n3��<��]{��e�~�y���m�x��A�.c��{�K�{`�2�
�a�RY%�N�IG$(Ԫ���\N����9ZP��B�V��F[t��vx�d�\���N�S)��C$��G�G��D�������7n�Ǻ�>wPC�W7Zu ���>
���k 'q˧}��@�	D�ēA��|�	�ֵ.��)�)s�Ig�=�|�4�$���q�UX��D���+�tM�����WF��{3zj��!��H�mCCV׏�ՀA��46e8�#�SW}l�}�q�I���"!rC�Z��]�h��� 
Y��1���i��e���܂�K���yO�,=�@����;n�b6�<c�R'a%"qR}n�U������^�����߻v�-`^�?v���y����c�S����,�?)"�p��q�����U-9L4.��	^�M�isf!g�<v[UK��b6@}�|�tua���o��-�y���r�"
����o>x�O!Z�E-��C �����|Cz-��_��e�>?�3�:񰈡]�o�NG�y�:�:4�8�1�_�E��@k�膚���T�<������C18N�h�o��"fQ'��,+��ns.;�1�Sƛ��v G.�N'>���r����gnST�Xh�	�̓�b8��5��,H�AM�wO%�&��Ti�rH�������I�^������Ǿ�쫠�����h��}p�A�ߚ`PA1��(��6��x���+�%1�����,8��b��~�Lh�L?.��)�!��n��\G�!�E=��#�� �+`�%��q���$�%5�+е���l�T���̵�4����MuhE���[�W�����߻���zѸgv��<�`q���K����V�)��!�)U�>+���dc7�����%]|����I�{py���lv��V/B$
~L�`dq7��%���=��qߤv����H���{�T�)�}G�ɠM�'��x�-�ʃdM���y�=�N�H9�T�tr���{-|zi���^�h���iշ{b|�*g���h�Ԙ<hR��c@��V����x�+�ud�R�n�\�؄&��ǯpC�����Es���gP[���� )�Z�2��@�b�^����#|�9Έ�Sf��GZ�u����*~�G9PfpK��D���W
��x�*Cw�h=��&�C��R��.m���=��d����|��,&6�m�v�DgL��*�z�
�6�Y<|���GL�N�t\�R�\"�fo�"-jW4�ϥO�b���TK��J�da"���2�R�k�X�7�US�5qвqp}��eʹЭ6j�B�dd:,�w#x��ꈚ�.�H�����d���q��D���I����_y:]�0v�š�/#�Hw�S�%�s������*�D���@i*�y�yxQ�Q��N9h<Ū��B�"��<��Jy^�	A��4.'�tzy�C�e���х�ÚZ �m{���.w@��A��[Ü���*�|lO+QRL)���[�'�$�,]��Dg�,�/�A�Gb 8@�--��۰�}�H�1}�7��#��}�VA@�Y�2����m�z��dDU]���q�5�6�a��=m��y�Mo֘�؃�5}>� �U�M=�Xg>��ш�d��P�3�W�[wL��|x@R�k�%s��y9�H�qWQĆ5(��\���P�ż�!#�4\�t��T`/�:r	��V�>�LY[���� ��7U*�:dmՄ����~����9UR��܎�dEQ��w����cz�k�����kE�$���K_Q�N�`(wE�#Y76�k�İO.gu�?�v�ׇw(��������=�j��{g�b�����*=׵{B�;��%-�uڼ��f��-;$K	�9�uZ�cfK��W�ǫ�@�h���]G�A\��0Dv��8�+e�3����Tl�fr��u�h�'����Ace�`�W(��0W`�E�-$�Qi�T�7!B�9Q�E8S�Zl�ml�Xz��\�xF���w�&�;'C��C�gl�D<���7��3I�)��NX�t͊�,��p~�tN�a�BR��\�~4`�;�ē�U�Zs}�h\,�������K���`��m�Ы�O����r����9��^���<�?<]�6�z�Ν�k�ÿ�С/C�v�w*���)��VO|͠��`x]ң�ǚ�}��	-p�\]\7^��*n�y�/���JI�I�=��D5��D/�#K���r�CI,���8r~���3�s�Q��U�v(ڈ���
 :�^ P��O�(���.M����Ȑ�)C#~7D�2�M�ˀ����S������[��GZ�0�c$���vsf��n"�An�����yEn|��j`J��~�:ʸ�!���nC|��AW|-�Eb����?���X����>#�P���Jr��ƮJ­,!�:�J���ξF���} �|%����<�͖��3̪�a�7^���oOPH3Ȇ��=W ��Xj���_��b%�9y�Fa~`����*�n�Y���R�^`;���M&�2P�9}�DI�]SNSk��X��Az��
��j�;���U�ZK��Q����MI	�]�}wh�K�D(���g�\UJO� �K�h�[�a�F�ޱ�5̄�(�a����6	y&�6�?�X<�v��6���i���6ȑ��l��.��(�O~�Àh�Xyw1�'n�����O��6�����­ѓ�K@��K�KI�F�-\�cl��s���h�ሖ�[��2ʪk�_���:e���+��9��R�."g�[R
�A1�uRRz�wL�Q�f�H�{�0�����*��ҩ�ҡ~YԚ!���]8j�Ո҈B�p��$��0Ų3�/Bv*��� P��C�m�j/��j�f�Z�J~�v*�ޡƎB���D>���w�W`�jw��=�^��X](���"�q��.�Y�|��ϰ���yǥ���Zp�F�s4����K�zN@yó>p"�����o�f訳{�W�ע(F�ޅ딧y�|ꉚ93��z��L��W>���}=��t�R���Q�g�K~M=>�*ر��|��[u7�$��\�m�)��XB'Y?���eZF!�XMPj	�-��Ⱦᅷ��}yLx���7"K$-跧`����㣐"�s򠷏bmQ��X�oƝᥙ��8��P�sX;����{U|Pnk���bQT}�XYp'��؅�����Ni앇�������Ө�BB���~V5;�!�^:�=sSԱ�":s4����%xӠ+��LSL8���P�D
`�[a"����q���#B �1����J�t}��s�n��9K�����\�Rh
�Mr�

�`����;h�u�D��x����c�LM�ǳh^vy����v�~M�& �\����@��
��#x��݃$�[�E4��Gj�������z�m\�_@
�ܮ��]�J-�^Ǯ���0+`�f��lW�x���� nI��?"y�x`�و�Ё�{�������W�/��`_Ak������9���s䵄}�|
���3L��^Bh|�=D�H��ja��)��鲚v�e�RP-EޏM�NJmfw�<�J�[���$�s/rF�!:��d~��S�7�_��1��C9��T����Mp�n|�wV�OMb�;��/���T��{Ɉo@]��m��ǘ�P(EhJ�t���E��� ���[���}��0���IAD��N�X�?�&|� YΝ>��@Q�<�)���YPq��,�6�V�iU�G:�H������'��)�m����`�r��uz`�с��*���φ�K�	��.�ո�":��l���<�1�IN,<Y�d�^��;��r�W1%C����lG�A���aՆ#fL�T�:f�Hi���%��ܕb*g_Nq�y�V@xK;y�BU�_��HӛV��܅ۂ�oX��x��Tn��l���'N�� 
��u�:����!
���<a%A��K�:3!I�K��3��!V�ފ�/ʷ�
�cG�m7��{��~����/f����;+�rCb�Ոn�����}�Q�T�0/�&��3ʹ>C)_X�����<m�]O�g-�EZLn��M�gn$�=(�Q* ���Pw\ݦ���:v�qmF�ɸӡhs�P2Y�p��?���Z�im^�&�3����75Z���*�b?h!��"܋'�M/�0�I��g�$?�X��}C���Ნ~�^S�S���b����5��������O��N�:f,p��WS=4�n��p��p<�X��O��ɉ(d�P���#��o��Ҹ4��=@�7L\�)���)u%�V��]B`Am�O�l��1��A���z�[�S<-����Bǿ�d"ܖk((3�ƪHC��-r��L�2LS�4�x������3�����L�:/*��^��!��9�ȿڡq���C;��o��R��yX���,t��a���տ�^�$Sm�w��AM>��t�T�1'7{ʍ�x5�_�d8ƍg9�����r���X^jEl�����w�~�h�	֠�q�
��0/t<��{�I].�fݏ�N����>?H�_�2~18v���3��D���W��Yg{��^�9��S�Ą���Uf�A&�H�:�+�~Ъ&�T��T:��k$D�jd�6�{H�C��K��s��&�j,��^�����%!�:W��6Ow�fץ�i�;�C^;� ���L�X��,�����7�C��"�MjO����GN��F��{G�\�D���t��Bc���������N:3�����{w�	�:����")��3�ͪ�'W�Tq�W	E̙�n��s�?��/�z���q�t2�a��3�8�����`n��4D�ʾ�#b!��7)07i_Ha�g?؂a�l���l������Cr��;F��7T1�[�Xn	\R:
�C~�j���e'uv�β?$�����e
�� ���fgN�k\���r�.f!�����b�+Y��ۡF�v�.U�~�0>���M�@!���VWM�A�؀l���*o��Zr�PN�.�1\����lwC�e�	W �>r�c�٨�C[seۭ���H�0�:xA{~�,�3e@��@����������S�B]\ R��Ŕq��Yʏ��O���Ȍ�$��3�Mm���V�@�E�@q2�@��'��7m�L��b�:����qĤ�$���㋷�X�ak'�����n+m��䮙����o�:�P�vu�7�u���%(���c��e����f��{��X�P�Iq��jᒩ&��h#3CNiI�P�.�~Dj�x0��Mk�e骗D�?)A���ۋ�����fQ=F�y%
��hZ�����FR|�ja�w~��A .�б�Qg����н�d�OBU�9��I�J�붥#��ԣh I���#n�Em�]C��5T�J������Ve���A͚[�  �-\�����K�)�zІܡ����F�ŧ�X:d��SD7?��:��D��%�p�Vg�y&����a� 0U���u6O�Y�<�O��]1�tiX�$��}P�f�IT`�5Fj����o�9a�p0&AZcp��'��!�IcOs�p�n9R�M�*3ؼa���G�*'iP=pJ��QJ�oz�~���� /��hr!��ʖ��Y�m�k�@vƭ�H⁥�K�R=E�mE�4�fB���q�$P06b�x��'}6ȸ��p�o8��$�q� k�;�IP��t�i؍'�lbW����ը�6�o�KVQ`���|�ȪD��*�����|K4n|�̽A�=����[8@�%�hӧ����iCN˴��H2�|\��#�NɢV��8�Ʉ2]ݫ}�v�Pݟ�qY��q�@���|�Οh��jj����%�5?bc�:�0�*���?f��V�wkc'��Q�\�Rx-����<�%�d6G��eƶ]f�pV�[@�̆N�$6�i*俑�2I>������fv}��.������ggw��]){ͰΚ^��P��̰��q�0��ѭ�?TXG�R�����Ҟ�3��n�}0#��)�2t\��э��3D��H��&�_�_�^3��IƝ���`�uf��a�g�" �f����:�5C��^(P��Wmxe��u����8��@a��U?�M:�5;��i1� �Y4F����x�g�R
�7��>��"��s�DƋ����X�i8g�[ơ�M5Ԙ�hL��,a#�1ܩ�F�q�:�)��6�a�f8�x��s�P�����$�vr�\-��@v�O=rTEw�Te!+����~ݧ
��G�Z ��L�Q�6�����e�UA�)�k�6.I8��a����\�<�����ܝk��ҹ<��J�i��=��{5C�����w oP�-���UN�<�l�s�Ek�Z�4�)tk��=s�
�m�.����_С4n���e}%jJ�O&N�!vk�M�t#D�[�OE-��x{]�ز��� ���z�L^�JE���+~ǀ2���ħǓ��^r�����Jn�;�"󓘚OZB^͉= �+b��BY�������(8��A�_����'9�.�B�r��(J#FۄR�6^;7k�@<�T���"¼ȵ��(��|�ȑ�.��7�Ӯ�C�����ߕ�']�RB:�'�U�hz}����E������l������=��F#5��s��{��(�I�%�44,��9�� ~?�?�il�{�\D���������eo��]�`�{^�$�7�\PY�ش?�)6?B�����|(@��q4�W��\-�Wt�]F��w
'mU�=�����@�#P�X�����RB��|Z��H�����A��D6�6-���\r���v�O�(��4���,������D���5B�\��s��6���d���T�7�j��WÒ�����FsU���}+S���}X%rv�,����Q+x� =�������q�s�7%�)���?��9�=��h�Y���&�DӋ�R1Y�A���< ��b��N�� N��������	���$�Լ�_��U��"���sھ0�k�o�f��ǽJiw[n�� w��*g�m�N}����.�:&�˦��Õ�)�����B��C�d'��.�uu?b.;L'V��t��Uz������K�O|�~��$@*�k2�􎿴v�*eDcG D�`p�|�a<�w�f�K��D_�L����y��s)L$�=�+��'�B��q���*��.5eI������H�	���ظ����<�'xY��x>�5`���E9:�}�0���y�<a"���B�Db�D�_����m��iC�����Ji�?�Л%�y�)�N�&7���ҍj��v~qo�(��ѣ`s��g#��t��V�T�&Н��e��!=(<��m�n����lH�j*���DWs�D�Cd��Q�i"���=�~�:��~��pH|�w�L���#��s��C"V��ֶ�מl��:��K��;���甏�s�����C�[��З��}G�������|���<��*	w�NX�4�'�]#ūa6�� �qr��Z���a��p� i��u�7�dqa��C�����⫂�.�\���١��:�w`ۀu`d�R���Eb��%I�aō���^���t�t8��k�&:��q�&J�q�\=�f�أ�p�9Ȯv� ����Z[/�������V���c�9���MSj%�`(y���5�+�O�qہ}��s��}ף��-S8�,����53L���,NW�#n�Y����[b"�e�'/�5�x�7�8�i1�,���:oJ����W�v,�a�K|~�<���HAzI]��+��Ѝe�a%qK�b��LlӜ́Qn^i>h� ��d��&s��U����B6��7L0�-ڌEu۷�\�|�K2GR��f�h�\���%�M0���Ui/d1c<��n�\�1��99),������P�_'���5�E��6���[����V�v�F`f��!�ST�S�S$	!�Mt����{t
#�z}�����9�x����"���I=3k��'��J�nfD�*� ��?������/5j�"e�cW+���
�>�K�Huܱ�gn{%۝��ڱ"���<�aI��ک���+Ԯ��p�t?
_f�s��^ 	wH�?4��=� �3Y~ks6n<��s��������t��Y�{\l�ۨ�.�d<���_tj#���Ϝ�=�|�����	�����>�H�'�a�O`�Y*4������n�nH���Yf�-��=:HB���y~P�.=�?�[��Q�$�4���W���n���uZ`��[`(l�m\q���Sp<C�6?�����f�&�bm1HV���!.t��Ê(ȑ�?W!=��#w*�)����|2��]S[�4����/�N�mq�4���!'B!`AgVʱq�w�؜����I����g�c5Q�~�s*��'��c;;�,�➼l�d���*�k��R	���DJ�ҧ�n �����=?F�6�bG�D=�8+�+��Z�lJ�j�[:�$)-��H���Ou�I�RVFu*��cF�|J�L��:�|��2�{�>��[�����∊Xu2��V�EPA�8��̩ݠ���#DY��5�RH��@�$iݎ�p�����I50அ驻$�@_� .��u�Ƹ��I�K'x��m���|A_�<�Z�#�O�;���+EE�q�ﴓQ�������9��	�uy�Йl����3�= !;�<�y�P��;T��W�L�G�l'������I�eӠ����@aLW>��F���O~��k�T��	�OS�(s�PL�|�hժ!ա���d����!�S"8"�7�ކ�q!���S���G�ȂBup�;��8��m3�5�f>g�3L;��-nx��Oq��d5���4)@#���qci�Zu��j7�3$Yj5�y�m�bA�c0���$��ߺp[-���8H�w�F�M�@3y�r~�^˛�ڙvW�ڑo�RQh��E�eg6������j����1خ�fX��ґ���o��u�[� C~�0��W��9V�ߵ��߻(5�f���!n�$z.�d�@�6I1챓R��jjd��o��(��ص¹?o��U���+��}���O.��~tQj��>>��(�����$W��Cs�x
�����7�3k�趭q8À맬4:�u�$j��bY�!�� (��&�1�T��8�Q�ir�B��VZ��U��i�6��Z��+��߲K���U>����{6�<��"�Ԇu�s4�Z��Ppz^E!���+����i�gO����u�<�תj��kI�ණV���"˘m��E����=�zmi��|!���O7IS���R�so6��;:8]��e��rV#M��5ޓ?����|�v�Co[>�|��ځ���g�[�\N穑�1��2qX��c-e]pf�ބp4 N �C����y7���;��Dos�x?{Ӻyq�3yG47,fU��0Vf��ҕ��I�
a������>��[!%�Ywur�Z���T�Mj�$�J�)R	.Ss��sg�\�Q�2��5Tʓ���QĻ(���P�� I>�Qf�a�P���c���+������;��J<�/��ߓdVo0H�s���k�g=���y����}�z�Βxw���I�B?I�T�|F��	�l�!�\X�2���e�K��@��\h4AbXDj�K�%��zzK�z��z��B�x�
�2�ƍ����M��ix�8F�||;u��+(R���_��E�p��5����������bY��Eo�G�t)g�8h�p�'BI�^T6c����ȘE����G~<�����;q��)�g�G��D�t�~�͸zT��Y�W@�G�3+�v�R*�*��ä́��]�p{|�T�|��+��p��$"e��kL�a�i���≨M�.��W]|eS���ї�}��.uW�@�æ�!&�k_�m]ح° u�V*(�p�&�G����.�[[r���D���\�}����c`b�чz����9D4E4���szB�	��hԤr+�W~F*%�P��z��S�K������eV���fK���Bߗ��w]v�P;*fR���)��]$@p�Ў�F����v�������1���p0�Sd����d*��!#��A��s���4��Z����Aev��Ng�9B��Q�_��x�m�f[k�%����d���XC��Ajn��d�=�����+Ĝ�+��u��9Fُb����s4n�R?��H
�0�J�#�ք��� }N֩%H�CK�(;�o�1Ot�NUEJ�|9�<��(��M;p쉜ǎ��Ї2��������μ�ˎj��,�  hN$�ﯛ�?��w�Rs���-�H�����Lh�r��`>R����b��7�8�4�����|φ�i	���=-��n�Oc`
xK:VD7���,��m�F��W��`W���Y)�'�
�t�n����˶�875f=�r�NR1�������w�<~��g�Iy����6ʈ��1��Qw���:�;2����緤V�2��tME�̰{�i�y�L����B��Pt���cLYc�9fa��peiv]4=�bh�;��L�%�%��l�Я��u�FO�����*��l���|���HI�Y��"���ti�m[I������.>�pY��3��#m3�x����Z�i�H���Q���b(�7�f�n<s���D��q��p���_b���=�[~�n�����*�JY��_���w���|q�4���g���'[��A�:�B�2x]^!!�]�z�ɉ,�Wi\�UooQ?(�,����ƻ���"00yO"ih�6+���q�Fo��5�7ũ�f���L8�9^���K�~k*j�	/5	8%���N]\����ާ� ���<0s	;�7B��-�����.�"���L���2����/~̓� �]�C�yG1���v�	▱��JR����g:o�o�+�;Z)�@��y�Z볖)?vs�#7��a�b2�P�c�KՈ����z�G�5Y��1�> ��mQ�`=]�����ѿÿ.Z���v3��[k����u�j^(�M�9�u%���MZ�ڻ��N㱛�f&�X�]7c���n2�������H��-ctХ��D3�@�g���R��cM2���p���!�E���&��H������VT����Tt�,���"�X��'	���86TO���,��q�����+eN�ӝ�2zn�g����3+��FA�t���k���a��)��$-�kj�={��S?��G�Rq�r6W},�m��&�i�,n ~�f�C�9��+?*�'Al�_5�H�By�>���W���%�5�?*���������ࢦe��Y����ೆ�iI���5
�-tfD�6hX�S��I��cm�+P,��,�*�C�&'����Y7ƭ��(}fFӈ+x����{�X�x�p�{��0�ix�B��H�%��W�i���n���8b ����W���"���54�jر�09n����dy]@�4�;J_+��e(���ɘ��:�Qъ����H8QK�+�Z"��F��bEO���3���ip�c6�g͢	.�UC< ��g� �>S��p&ԕ �h�z�U�����U�����Cm���S4j;z��/�:�~��h��n�f��L�4����:��~�x�A긲������=ya���Hg�Xa����xŢ�����մ	n@�e4~�ӟ����
�ag�X��sK�i���Z���J_�+����O�G� �1@��jt�J� 0�� ���E��Qߊ��	�KHͪ�s�?Jt{��Y��g�T|��$��lm�[ҹ�B�r3e�������3�6�V�� ��(���%:ˏ}*yx+���x� �h����eI�)��V�k�K ����M����������0 �$���{R�Ȅ]v�l�D3a�l�j	c�a*h�F*A.Co�K�
$���L�������{�5�j�}[6��~:Z��W� �ӜM�|�3�������d�#�:�7'�n��q�9�@�E�ι9��8?����Z�'�ό���r�M�b"�]�)xX�c�$�5�.5hq;����f�xgH����J]a�w�j� %i��y�M[hvN4�&P��9:e�ەՋtGU��bSQ$f��~�!�(߹������8H��#D�������[,X���<ĵ��)�ŗ�/���/�����͞�Us����O�2ӽb�t��;M��w�	�s�T�M'�sG{�`z]�G���&K��x�E��B:V���="�k��+�[����^Q��<y�ʓߐ7���>��2`���^{1��
B�v�h�&K�Z�]a�Qu�\Y�瀰K朞���wҰ�%>&���0��4	e��%�l��=cp`;�����[epP�����LL�=�Y#*
5�E�E:1�JN zr�Z����9���Y�Gh�ܤi7�������5�hF�m������^.���{���DB�LR�Y�_�wW@�\7�n��@��s��'%ӝq/w�������l��:H
�u���=
�HZm���K!�'��vy�-��귬��)
��7�`�3[ĜD/Z���!�B�Kz�|�j6	ZX	.v���#*{+��KU�����G�����B�%�㌶k��bFtҙʨԝ�H�d_��wǋ��_��6oR����ȸ"����ARݒૄ����};�C7�W�la����4�òCr��̘q�S�@'��b:z�_	�
C�MqvfsM�t{K����ςk�z@+�`&+
 ���Ʊ,��k�9%��9<�����5��۱p��HL�#�O8\H�B�b�3��nkIj�,��{l����3��ݞ7E����u�*-yMު�9�[N6�]���*ԝi	��6�-۷����������Zl؅S�������T�E�^Zoh�(���q[�����C�% �� #!BKO$��JI���i���\�<�ԋ�J�8��n�X;�ɗ�e�݈q�CI\m��ۈ+��7}�N �K.K�s��A��9#@Ë�|�m	o'#��G�]-��W5�L��[M��!EJA��ƪ�9��G5�2�xR�^��q���xQ�X��z��vaTV,�O���Rȕ��gu��>u?@p
��%��Aׄ�����]��r��#�&K��d�7*߉��Y��J{S���:�iK�!���BeƸ=e1�l�M1�Z:A���x�H\����V�\�� ���;�JΊ[ˏ%	��	��fY���]ɭ�D�q��}��+�}�M@���qꧢ��t8��m�P� s��:����:=Ya�d��;�_Q���k�����)D�8F޿��+1�I�\�ڇI�Y����i��)��Q��kh�.܂��׎
���!.�v7R*Z:&�l����/���w��h�e$��*�H���b��1�0��ě\����v���(u/�u��B�ऴ_�΢�3��B.)�Kw{%�3�m61�?�ZL��M\:j���%�k��֘GDt�����
�P���k�]E�ట�Ws���E&��	)N
�4�gq�ߟ�����5`�Y7Tɼ��M.�4�9�R�{e��j;pS��~�_�j:�������&��#�t~W�"�1أB9���ܧ�ߏ��zp*Ǡܞz�!�
p��9��'%������dlv��"ýfw&\���A�J㤟�:!��5�����t9�
: lAY,�*�g-��AzU.~���#9������5����Gs�x@��%_�7C�U~'���0�"�yY9�
��D+����-�Xۓ	�<K���\vs�[���l�V�{�Q��2\���;���x���s϶���令�k2�$�N��.���p�]�#i,�6[XZ/P��K����Db��i;a2�z�-���Tu�y$klg�>�[�V�?Bi�0���Sa�oL�kpmU�����u��H��Q�h݋���B��Y�ؔW��fL߇��i7���@��u2om���. ᜘��ᅕy��Н�����(����.3W0�����"�T��e�K�����aT��?�I�#^K56_d�[��Q8�R9��)���@G����Mb� })!���w��'�ٰ6Uv��+�rKF�2�t[���rd�/�K+p�Fa���~�9�8�	[��-�ԧ!�Cy!�Aਁ+�È�1��AAUF��Kҥ��7���1b��*�����!�,��Drp�ҧ?@��]�;��yG|d�6����SH�V��=��h�wC����{�Wv�w�u�(}�J���mIk� @)A��!y��Nsxs)��=�d���|��b�+k����b�@A���e1>�c�3b뗩��@joKt��U�xHmw�b1�0�d�%��Ą�Mxy����F��%����$v�Z��2��ȿ���G�ߠh��;k�ʓ����8/�&7�@�
f�%�?V��j�hL�����~��d��x!!���J6mmM�a���Au�$R<#ԫRu5j1O7oҌ�X�����MM���J�W:�BR���B"�o�Ku��--_(�n����S��ŭ��6d�����ٳ���X�?���>�!j�� MD��c�\�4y}��i7(h*<���i2��:o-q�ݱFj&[�-OY&�7=t���@hقj�Y�~�0����G�=3��v�e�c������i,��R����(^y\�eC#N5���Ph�
<�nb8[�π6���L谄���6������-�x~��J����u�I���X���h�p�KK��ۆ��&2��pڱ{oI�����*ܣ�Р >G�)�w�Z=����Ϫ�������,�����~<큙#��r�@����
I�A�t��gS+���.a�HqoP�v�3��qxL�M���e����i'����m;���V����H��uڒ�ݺ�u!�������J"�ە����9�{j(��2�l�c�0�)��I[6d���u;��W��w���$�?G�����w%����Ùs�N�5�����%!}\�����TJ2�â�#?aQ7�v�yaC��%�䛕�r����7h������q���}P�҈���P�=�O�:a�n�)��F*�w#�LC��v~��Lv���ޑ-�Sd��w�Wl+�lZk��/��(Tc�>2*��=�F�﷽fVi�%ZO/���r|�,l�?>0�?��<���"n6��>�o�b�.ņ"v}����=�7����H/���tI����`�72��b3��R_8Ë*�y�%�jvR��U�q�@Ӏ�;�B\�*�Ub{q�'�����J�Z����PG�?�"׫,�@_�i�bI�_Ȁ�I��a|$�64��@vp>mxA���\����V9)�^�U��"�"`S���TV�iuĚ�r�$���l
���A��c��5��e���r!8�a����<^����tO���w~�	
���b��s��x�ā�1��jP�B ��Z[�~� ?Z0�ݓ5O��|�l2�i3���^�l����+�����lIS�����E�դ%ܤ��\�ܬ���2I�U(t� o�Pn~�b2-T��9n����c��3�wq�v�mU�93s����!�;��H�����.T�>L������'��E6�ē�%�Y�]lZ��N8�>�����([�ֵ]��p;�Q!	���Pk_Z�@����N���#�A�5����(��{�"��z��о)�[,��p+��(�׀4�x���֛ϛa���K�@.DL b}f<q(+"?�Q�[�Z�a�������O��xg(y,�U{�7w���������FE���"��?l��2��4Az5��C8�+��V��U8N|[�:�M�%m]���JUV֯�?���+е�����䖀1&��*��I`1~[�z��x��$����JB���Q�=��qel� �t��9
�Yҷ%Qe�HG�fI�k_���7�{�L?8�N �!���t��~)}�����ۀu���B�>�4r@' ����dav��I��ݪ��:���{���_~F Ŏm��y`b��@�p2��bO�Β�ԝL=�"�]��%�c��DÕgB�9����?I�݂�k����p��bVO,�ܓ�)8�&���hWg�>�ϭ<���_{с�0��|-�e��I������ܑf����FA�J]�
�����9�J=c�4/�@����؍�רI�umخ;�O\���;�Ue_9������X|�:_���5<���Y��V:�_�N���ڢ���O��>�!�{V�-,5y?�N{�㌕�`.�S��],$%/-t{Y8e ����4�`�����{K㈿-o��'vv@K�R�|��޲X�l|���~���;����9mb�$��ͮ�-OT����:�I��yX�9%�>�4�N�fI�Z�[9�𐧬��&qe���L{U^���,�4��\�!�Y2�������j�"(��F��U{��\�? A�V��?
�����	n�oY�
�u�%SB% 1g��Y���I&ðjl M�4�^��N{wJU����қ�TG��C��|���@n�ٳ�k����,����kK��ۯ�Q���X9�9(�zID�('�:�dD� L� ��a��z�:�}��V �>�|2����GӕtZ6#�t
�m�_���W��`��Ɍz�8!����;���;�X�~��������i�W�HjW��,Q�����+qhzq��P�?奖(J�=���L�����n���a���J�cj�Eb�
Q���G�e���$�K�_O�t׎	P'0Ð-}�NS��Td���_MՕi4<�5�Icg?��UGt���2�E(NP\/*�Y���ia��'R�er�B�+���x4��_��Ym��P��1���8��Σ�y�59�XࡕL�)%��%��aߨ����V-�>~	i!�`osmq�</�����	H!'T��7������ɉ6�c����Ρ��}	�x�T�B��Ƀqm4�T����a�qf����8+�yG#���צ�.L}��֌h�;�pO�?�S�7�ǧ
���y9u��C?Vs��S�$s&��b��e����N�I������|+!(�&q���$��?ɏ���~��O�7���G�+��L-�dH`aO2��jH�_���l����!��������\�{kW|�h��F^�W�*f��@<o��TRJS|`W��^K�s8D1䧣��g�e�D�5X㌲�CG���;uaO,�Ω���-`s��C�e��1f�oUavk���!���]w[��蟆��k�+�/����|��ݓ���9mY��є�(&�D�k�ͭ�[���ϑ�������ۯWN��4�U�w�c��)t}M#(<�~7�(���˛
�ó��[T��?l�<ƧeѻK�,��3��lk,��<F�
��k���U�A�]E�;^����һ>����sUU!��B;k��&Sy[U%] ����+���X̠z��=�����@y��&��<H�ԁsG�7����S�Z�P��&�|�:幃�/���K����p�����'<�0='
�)�� �,�A���]�ʮXA��~��R
��պn�$�C%�Ц���LU��'��M#í�ϒ�_�F�#��\�%�4���"BE Q��B@,�[�SDi	�u�x����M&]��M���<P��v� ����7 OVG��!ls�
@����='���c��ϴ��VU�4�!��S�(b����/j��D~�\�-wX��	!Ӫ]Y�ކFS��?�@�QU��+�3{<�A$�Z5?#+�]�+i�AĦT���H6��~Et�v߀�j��q���O������$n�󥶾�����<�lj��Ǫ���q�y�{�J�ȦNzR�agC]�H�񵛎r}�/	"��[����1�>�k���qM��Mq?��vtQ�	�x��gƸ388������|4F&K���-Pcʲ���Jƀ���cU6R�̖�d�F�D��'�왣ץ�tu�o�!}��veoa��Wt�K�9�x$�L;�����p�
#�	�,����nD̚�,$cٙ�c����e�l%\Ş�p<W[���<@�c)h�݋7g;��ٻ�ީ�Z� H/J�r�J��BQ�d�$ 
���GMr�B��$��1����p�s����Q\tɕ��ѱ��Hl-
�'�_bJ���Oh@���$T��W�͝�67���<��8�6��g��K��/v���ZKȽ��!�����207+���1�.����p�x�I��`P3��t�؎�%NH X���mˍs���D��oP������<Ba�sg7� �v:�f�M��Q���!����s��F�e%�U8�;��M��n�䏰Bm�O��eD��2����^~Z-���,r D�6xN��)�?�POq54a+p��W1������W�5�N���kh��]�SOwp����C�a@�u�<Tg;���-`�jF-�pF<B?��Q�PZ����Jlg=��-AxSy���p�Vp0ٓ���Hr7<�?�,M�sZ�@kk��w�T��6���}04uwp@6�t4|�ƪ4��:+z���ے� �t.u�_�ݍ �UqB��<M���!ץR�█<�c\���o�;�@�3 ��
(A�=�^����Bs��?ʔ�.�]c�����X�Sc�+�LB�����M)�OE�kL�եW�u�U��y�s���C¹0�J��˗�p�D�Z�p@�d\qfk��	�l-��%`�6��a:�o6x��j]��*�����O�?��M�8)$���8<�g�b�:q�P(��dO�WDN��c�p�n�(����v��I夨����ܦ!���Ĩ�E_���'�u��"�qH�?H�7��/3)�D��J�e�i���'�D|��M8�3a�?v����60�o�PĆ�Ev���>q�zC9\o�ʾ((O�v6�5 1A`C��6C��$P�x(� E
�qRU�C5�W-
��΋5�J�T�|r4�g��)vE���Kx֣�L"���&0���e�\�ù��;��)n�<	��)$��a�|
����.�d���̓����,�E���Y���{���H-#�V��(�.��ǑX"�t}�b.O�.�m	K�SEq�֞�A(�Y�Y3ٴ��`Ӎ�_�祣���|�9�6K���C)��d�6!�<qOC9���\�X!)�l[�A�N˒�*2�nkgx�)�׃1S�vO~�w���}�`3^8Bg�F�<7������z1�Ԝ�s��	�q�
s���Y������[����0q�ݬ�?,���DB�4mq����\���)�x_?ت���ZU�V��x|��B&�)�l�"~�]y���:,R����_��I$�_#���#�{F �0t��|�!��aR9ф{�g�򻢜~�[��(0'`��I�I�5I���X���_��Q�~�G�W��A��D�t���S��O#wuj*��3ܶ��U�}�ڋd�Y��,O�cS�,���ML��%i^��DV2��ُ�MűW.c�D�2m�/B��o�mZ�axh�Z��?��eY�X��_1)`�X��eq
���"�C��Eb,]��#o� �v�F&R�8��o�q��:\K7\#4�C����\>���g��t��?F�P�(bO���:��u9���30�E4:ckzj�BO��x_aok�t6o ���:m��`W<��K�hH�L|��,ket�m3ſZ!p/�L&l����s)�P�8�o�c��b>�������D�Ft�F�F����	���,5�����~L����Ӊx�u�I�(C�kܙ9,?,
�
לF��`�o��%f���1��5��Mt�0w�M<���vyѢ�Cπ�$�J{��\@O8L2���^%�.gf�j�7W���t�K�{���Y��|�Se���zT<:����M~�+k�*E�L���4ɢf
��>G�E|�{Zu�hr,�Aek;��� XOL����&��l	�E:x9��G N������j�K��̤6"=�FTX��!�coLh'<�
K
$$@��P�Q��F�ɐor*���-Bf�'���]aa��EV�T:M��Cfˬ���ex#����a_�[�S���m���G1��U�7���(�
Q�υZa�l�=�{Q���A����ᓬѫ��#��W�\} �ssI�g�J4+!�̟3�D�A(�+(G�WE�ϔgE�*�M�Y��̬3��i\D�NNߊf��1y�r)���S���M�;᧟h�8Fk�5��">�����lq�d~l)�2Fך�Hu�w�NBd�W�����_����.�QFq�&y8'��xn.0�S�\7��N�$�s[�U�e+�[��������#v@����.7���.�^��c�T�pc ���
 �{��]�%2�OeJ�i���"�Z"��D�����lV×^�l���@���o�uoҥ�SzT�o�k���%�x��݌&<JlOZp�ΛGa��t��Hړ:�r�9du�����u'bl���<�ʥ�,LrX�[����$����i2uQ�SFo�#���OtXQ�I[��	�(n�? ����;y�./FU���M�UUY%q�[	gEJ�{�>�5��{Pf���z͢�r0�kA	��}7�]�o~���t�c�s��D�i��G`��-�r)A��:��0�_��T��9�
���?j�_�+e%��8Ǒ��Mr(���t"�2��8?E=���댳5��*���	2I�PF�gf �D_�z`He��#Z���1׻ğ��"a�r՗�����<��A�@]h�D�ۓ{�?�v:�}�r�� ���0{(� ԟY��G�-u�J�^�����9[���T�U�Wt� ��H�/�p�"�h�CH��x�|F,���^�B�<آ�X��s�y"H ��>��	�X�N�`8y�� J����"���P�M�.��3�hUa��Y\�,���/��8����F8T�,�Ct�>����������\�D��i!8e}��i7�y|B��Ҵ�~�9e�͔s|���1��l�ÿp�������i�b)`&D節T3���!r�&8���*���g�K��$��@�T��]���s��N���; ����9��x{� 5F�cbP_%�c��[t����R�Ѭ��>$�1�D�>mt}��&.O��+������)H�6�3�H�bWH̀Qhʣ���Q��C/_%חA膗��'��w4[�6>��`u���ѱM���r�u|��@v`����&N�2ʇ��0ls�8^����w�??��[pTv�����kz��u��;ܓ	A0�*Bi�O�n�T(�j��'��o��pW�'oM��V�\�Pyq,�E��lC�����R��K{3�h�z�����,�A&-Nts��Z��?^��~V�$��������{�5��+�X��
��GE���� 6�Iԉ���?�>������H�k��t3�� ���.�ls�JIL!Mg�9츶bUtP�nVbjՑ5t������9PXA��ς4��P�r)�M�rk��Χ£XXZ�Tr˒����䤈)���3}����X�jej��<Ra,�P->]�;8�w���B��"�]���e��=��3�F��J���2�����$լ5_���Tx���`Z���&���yVZ!������(M5�O+��+�(h:��ko�/�*+lJm�3���a�(�����"�*�t�D�D�%o�4D�¥l��?��d��?g��#P�7� &5$����.�/�ua|?I&�/y����-�Aw��85���XQ/��]r���/k�U��	5�U�����]�5B}]m�����k!C��R�^��v�F�YbX��_�J��_�Ȋ�XS+��=�;������#�S1j�GZĂ(�,���5KS!�M����P>��A�ik4�@+��5]��&�	�V4�t��5T��( ۴FUYyDF�����8�(b9S3��Č��C��I���$�b�(��7㞀eNx֎��~5n�^Ꝗ� 3�=�%�I��;hh��5�����o8�2�G�v9s��9\�d�N��y3��(�����Qh�>�tZ;�W��)H��a��P��K��\������oU�Y+�����'�3��������Gc%�k��و�TBU~�SU���PGsUpA��[/Z����m�D	5y�S�R`b{s��y�b��������y�N'ѯ��1�1�7����8��
�������� ���F4��B��D:T�%�����YKZ��J��U:�(�M��~B~�+��x?��1��IOm�����)�I^롊�-#P)�����.%��ދ�h��sT	1���Y� f����}!BY*o������V������9y�Bs��F憩rΧ�^��@h��l����?_S5���z��Ī�ɬ"���I�$iŝ�N�1�z�R�څ�x�X�`7��9����l�7����b��������RH&g�ƫ	���h�Ĵ���d��*�w�1X���]���,ɑ��'R���/�hM�R���xB�����0rţ��:N��O�jV���y�d��~/ѸG�ά'�&3�sQ-�&�{�͸�s>3`\"y㝚�(�ݹv��w�x!#�;ºw�@���.��>H����0�*Iuҷ��8װ�(��U2��={=#�M���҈b��P5ÑPj���'ٻѮ�4���$t���ĩM��{��K�Xw�J?��a�r�4�-Iצ4�"��|������Vg�VΏ{��ߋ��i��+X�5q�FwO�k>����?vw�� �XY�f�+8 �i��&q���]����x��A����cWQ�2��i�h��U� ��~�yn}����/������`���ҭ볔j�:�\#���N҂�M�Q���s:�Hp��2īb�JǑ�i���1� �ƈhs3�]�l����1fq��`/�ޒ�j�V�A�Q�����ϟu+�6���5V�!5��o2q����<�y=�����V;�X[�B
*��e��λa= N�k��+�^v�4�v� ,!���~/�(�YO�?�����Hˇ��}g��q���{e��L����ll)Ԃ�A��o߲�C
(l�ܜ�s���
�i�g2c�ED;i���w���שf2��>q5t��v�!&;��)A�z1�B��K�#L�5�{Jz1���]����8� o`��?L҄i�\%Y=c��A:\Xk��D�|`�����t������\�V=9F�l���$����y)p�>��	�T��b���[C�ę���sMM<^��χ�������eSl``�� �;
�"�fH�6��/{�|lc��db���� �	@涔��l|���3͕7{2�o H�4w&'S����7���,�>�Е�e���E���s�2�����_����\�.<|hA�a����L��.:K��>�6��r���YQ&,v���E����]@��L@>����KIߥ�m��G���:\�c+�	�7܃�Z�<�ep[ڄ�����YA��.X���I�ƓQ����SnyY_����'�F��c�������'��0G��ޜ�-F���8i_&���d��i�An
�>M��D�����C����*�㘁����i*t�G�
����[���#5d�������ԪA��",�6��"��œ뙔�T��kw?�M֑2g;�H�=��eB�ADڄC5+@��@rz>�J��GP�>��U���p:h�yǔwm�y7��ɼ��l��+Հ`����H��*�먪ٽ7e*������	��IDC���!]DR)�!eH��Շ�JZ��O���dJE�u��+��1��'Xυ�6T�X|��*�uٜ
�" �t
5U�d�/?(��L���F�j�!��.�׌��-��|C�}<�MJ��O�R���8��j���n�/�w��`��6gjvr���OIG�˥����um����!�>MPW����R��'�=�E���Xg�@���&�;���NW�[b�<���W�L~/I-w%�0�Ѷ*B0��';@���6 �.�b2E�o�ԑ.s�������T� |I�1��)�*<��󊷜�b!�P���l�NW�_� �ջ�m�Q'���6E[T�t?���I;�����o˫�h|#���T����r�?I�)|���G����+�ʶ��l� /""��D�OɖLn�TB.~
⋇h�L!5�r�sTo�x�O��E�w{�#^YiaRZ���÷����X��f'��Cܫ,pJ�s�C\�}[����Ց.[�O1���8����Y��l����nR���t�`�ړm��հ�u������۽�6��{+�л�7�~����G9��3vu����/Q���.���%>>5�ԭ��.sE���'/��ʄK34���V
gh�b䩙���Z)C���Pk��P	b�I]_�N3������A��"Z������)8(K���>�������,t��U�'�ΘB||
_�����"*#�������k��U6��
�A�߆5�`��TH��j�Gi�8�ώ:�j<�VWpE^� ��k I��I7�J�0�wa�^��tH�ڐ��y��� ��άs(ʂ�e�C�pC:�vzB*��֘� c\�@z���Ib��wSP:ψN�-�v4�|]ڴ�Ҿ�\:�U�|���� ��;`<�R{V*��#=T��J�u���S/_	1��mܒ;Z�1�T!��F#i>�%�r*&��(��)h��s�C Ab���_����Whʫ���t��Ҩ.D����ܓ K������*{д�>IL�zQpzͮ��XXF�C��4 ��86C�ܴ ��߈5�Z3x|Ng7�
�kA��,���#W+�QW��k�éD0�KVSq�0[P"Z9}��)�,_�ґ��ϴ�iW�;��!|������1��z��	�N)Y��4.HJ�1d�Qhy
 �_ߴ��v+q��vLc$#�N�r�_�5�d����<	>���Gx�F�'�hOX`~֖}����-�Ի8�D�
�����IK���~�}T��2�S!�r��r�Df3G�`i�E?"|]h�{�����Vt���Ysr������.���{�)��~!�K�N��Nï~mǪ?�L�_%~�ɑ �Z ��"t&n��k<Pd��Ʃӵ3�*nI��w�|k(�i�O�G�6��wؚg�'��z�hp}��R�8s�=7kv�S� N���q��	�D2~�{٫�m#/�d#�4��2
�\�DyCz!�k���X4<�|T��/I���{�T)�!Vp��̉��|tCf���I��
��#����:s��ʰ����1e+�0�Jm�;���>��q�˔L<��"vm`[$e�<�邦^��Y��*7��t<�-t,�_� �-��W�U�-f��MOkfJ��@\S+K���.�/�	�UL�تF~�O�����(oWX�����V����A�HZ�P}�(u7T�5���=��7t	��1���X>��xŇ:��|�0�^�MÓ́S������3��s:Օ@�C���� ��+8���s#�W��b�f$��C �����W����/$w��_�x:��E��X".��b���v��2�W�L��D�U�Ck��m�胰����a��+���T�����(�kH4��ȶ���O�FS�Ʊi���+�Q\�i�_2|��Gȕ�F�O�;�]iغF����Kc7�Ύ�)��4j�?��F��.Y1(�����(���ꥬy�KF5�H�bI�+s��R$Ŭ�"��|�N4D��VX,bd��"9�]�L���w�:��������M�l;��\r�)�D���l�/:"7����u���H�q�wBW�a"��;6������CqMQ�H�n��#a���|�9r�x�?FR�?���Y�ư��-��3�q���Ӆ�}F�
1�����S�ǭGL�Eq�gy�<j���d�R� ��*jA˾��NH��]Pk%��W�N1��<j�����nχ����o��T�̑$�̉�����T&�w7��E����̀�6 ���:��Ut:�jF߉�j�s<�l��|^,�LG��=�O�׷nb��k��^.�f����y� n5�8B�|��"����2縹��]�����G��>�?��n�4Ie�mFA6[c�e�4&�����t�PFl+IGo��-ްW(�{�V4��v�U�@.�|?��6�U�;a]�'E����o}k�8f��	�"?p��8�\�$� `��0����_��d������`��\�9�[J𻴬I�=܉07z���n�������dQu��:��j�n���z����_f�����Ĥ�^M��K@�� x��v�uN���z��N�w��G���T��ٸ��hY�IZ��ؖn%e,_��,@bq%��Uy-d�
�I.�ʏUD/�D.*������5��k�`q�<<4@�0eqT<��Y+s2��t���}�T�iC[[���.R�[��
�EQ�KϏ����B˕Yv�M���I���QK���������ܯD�É�+1�d�*c^FN�]C	Ha ���JO�n�.���7/�����ЭG7̲�A�#����dj?0���"]� �`����sw��{�Fq�n��2���X������R����cXM4ڗ!`>�-�^�i⮰��]|�SE�ZŇ���%L8�3�0��f��.c�Rb��=��'��G�ΰ�y^>��r���t�8�Rp�]Y�4���Ȼ�C"�0$86'ao�����^t�'� +\��;T�]?c@1�bx�U`r[����'Zj��P�1�9xj ���h6dg���\\�*[@���D������*�o��P��F�Gh�2+���@]���C4�桝�� �"�hIJ7p�U�b���&�3dQ(����c�&�X�"L.R�e��I�J�&�����`��eH��8�5��ߢDm�a}��w-B�r��/2�(�u3,�!z���3XB��Z�VkN,W���Km�Me�T����F��±��Z����l��SGTD�4�Dk�go�<�S挴 ������ʢ��M�SJH7� �9��ҞM��u< �n��{ܥ�s�D�����#䛇Rl�H��,^;Ҟ���l�
|��<}v�Jh&M,���!��w;n��"A죲�#1�Sk�%�Q<�A*A2C3�>6���붎k���Dm�f�W�s��\����/A�n:�ʃ�m���JBɡ���D�Ͼ���0 �f�I��lM�4ō���3�l>D3�X�����6DA]oUk����(y��kZZ#7�c����K���ġi����y�f��?Ǎ,�h��+d���Ӳ��M�-=V����g?�+��D��J��FOh@��m�\�J�p�g�˔��7ay���DO��I�}Ƒu�o�6�7�F� ��z����r~ݟ>��N���KJ�!s��艹�$��*�!��q��i�� f�R:���WR�q<A�il%�������X���`t��Zf~�V�^^�����ɍz�2"&��̪<71��cܷ�C6{N�7�e�������I.��r� }��ow�)�� ��#�I���L�>f���׺{4��e��,4��E݋�?t�:h���fhM&��D��{����*�52���9Glzo��]�v�~Ѥr?�v7��%��a���zZ�H��ҷ(�|OzH��lsH�� =p6�΁�_���=�@׫�ft�In��*{�&�;C7��޳��{^����nv^�0�੓Է��uCN����-ޮK�'r�S~����y�I4�Ij�=c�K�3��r�k��%)M��L��n�$�CQ�Œ�̑5㞺uWDsi��ڳf��ݑ�$El�����e�&��H�I��yWw����6`L~�-Q�T�1O�N{����y������K��|P�:x�[[��Y��c���U��|F�NZ��_�.�˲]�;b�-���q�N�-8�>B��}�dx`���(�0_�?��"r��X�	�$�p�w>"45��;)q����QZ;��lLw~ ���g��қ�[���-=%����D?S�ׁq�㆙#4��v�vl�K_aK�y8�th�%�O�D4D���}Q���,���)�QD=Ez0q^Y���Z����bX �ʭ7�`�����0�\4���ԯEe,C48�l^:��R]������^R�α>��C�P�n�Y16P�G �NQ�L˵=i�Ih&̶���ˇn%k�
�ߥ-��"~�
��P�(>X?x�OJ5"�Ɔ�՚5�p5?������x�4趼�V�b	fu��o�{�5o*�DC,���x�8���@)�iO9xk/NOZf�ƫkNF�(���A�H�d�"~b�*Vi��K푎�G/�3a��gs�i���vb0�55M3�]S��ӧ"J���Y(h�7z�/��:�R����@��_��%�4�yQ1�8���	\��gj7���熵�jP���1�����
��޵���X?|&�tٺ͑_�5�:8��y�h!-P�F�����6�%�%����%y�.�9���?ؤ����>��_��47}5����G>Ֆ����h�h�kMp�^U�b�<��(2�­��Nw�9�y
W��g�:��;�x�^���Xq�������⸺ڗaI��$܉]�u7֣������"q�Ԕ��8P�$�+9�@y��#,��z����g�]��J�l��q�8�.�D��潩���W���I/��2�I�[�I��@�ny�7���YQ�]�i�u�i��)����f��z�u,�.֔=]�'k/�7#��SL�S��K3�brx���
h����A�L����*�<�0:Y�8Ѡ�8�)��q�4���u�B�|L�'fp�ч�]��������C?0�j#mx�uP�4�w��YE�t8�G�;��9�����B�����ŭ'(i�y�N�����}=�OE��	=�"��9�(��U8���4�e�5��=���
���%�[��B���8��3&V;F���Z*i'�h���
-gD}�+z��D��L���îZ��w��X�#����C\�����7��dsO�Z��r|�H���p�`	���#gC��Ya8��F�]�C7�8�/O3dU�ɇ0^�k��q�/���i[4f/=�p/`T=�C�V�F�ZnEAg���IoNW�����g��C�����R��Z�~�0�����Af��Ğk��JL[aG>qd�Yc��w|��P��Tn=6���?��=�E�5e:��5�ȩ�:��͂aW��}�lW�A����G佬�'�>
H��J�y��8�0�I 1`�P�K�����6�⻾j����g�)�9��p~:�(��w�{j�B�@8�	}���w��,<��&ő-R�P7]ҩFy��R�!�mnJ3������s"�Ҝ�A��>ϗ�D�z�Qm�x��Kø�B����[y�He/�!;��][Gʼy�z����mO�L�D�.��!/%�(Ъ����iݗJ�b�a�'ut�G��ʢS߀�� |YJ%����Wcg��D���TF.��[��ga�Q��k��w�_7�ѫOyXGc���<�[c�]�����>�>g������q�,`C��ҥ��7[��,���Y/��:q�0v �� �6z���I��a >b�զ=Ě���QȲ¡��ܧ](�|�3j���{����Ug��<�x�
�_�m��V����WL ��#&+���$����3�0[�3���\C�w4O�&H����i���Ko�H�n˅�pB�KT��w�#G����ـ?ź�ڗg2dp�m���׳��!�X��L�����c�Or|�$�jD�o��{֑'f�l$�^?��Mi�Q�(�dK���jC�.�Ɔ�x[ �N\���}NW�,E��1�YX��7!�QP��dۻR� �e'4�d�B���ǀC��MU;j�'��t��la���ϲԄ��Ⱦ�����0���M��1C���8ShU��$<<�%I;hS{�%1�Fu��o��,o��;i�2y7K��>F��3w�"{�a�3�_�+K�2Ie�i�Ci���߃���b26���|.��K���re6�q$~�ȑcً[��EZ~m���t��_�;/)r�t�\�Bt����<5(�
���jo �R�������<�F����{k��<bQ̞�Z�KkO�i�S��FTHf�gb�'t�9�	$���F�p߇�5�5��WI��!�y��a6EǬ@xt�z��p�I�Z[I�%�YnF�PT�0tAy��As.��`��T��9GCG_�,~ ��n'��t�ƅoa�??˖\(���ʜ	P��M�a��K��:l3�_X�e-�P�4 ��1�k=�����3,n��3U�'w�g̴��o����A�{�j�l�):��v��J,�Z���.�>҂�z��|D0�*�3����p�0R*TH8�FF��O�������6>j��0��Y��^O��:,�A��M��u����+�owN2;�%��� ��$��]�Z���Ţ,@続B�̡d�����:	j��~�i�b6�$�L��A��K;Aj�؏�j�Hʔ��j�5�Ƣ�LR��3����^xųx9y 5=ۼ!3Ge�`�Z�X���L���iE/z�ׄ�����Г��_��8�Vh��fPݹ��JŅY.xq��M'm�j��5�����4"t���
�t�ZA_*�C&_�X�~�J�?���q�O. m#��Դg *�^�L#�eY�w���M�"Ӣl{e����zy+�S�>1�Z .�I����>dJ�˵�T���>Ds�9$LEkQ3F[]{���N�;��8���� c,8�A���qT����>I"�'��l,����hgIv e�U�T�p�Y��ԥ#Ŧ#t���#Zh�*I��!,�z�ˀ��˩X��ҷ�I��.u���1e Z��J�.M;�[<�W����0){T��Nz�����iZ�?���>�R�U���w�8��𝁧��Ȁ��z�"�'��{(�,ZC�x7<`9��G�g�
����A�����#AKY�:m1XT�[C�**�AH�~}�X^�i&�W�]�����F�^�h����v��ِO�}��mv�.����Z��~��B�w2�\S�����>V����ٷZB~�~��U����i�"c`a��J;<�^?:�D)�~��|ܕ|#ܐ��Q-d���P!�X�=�b��k��;E�&���wf���:=���Z���bȣ� <jYZ�����*�޿?�	��V-�84b��L����M�W�Z[��%�Y�;��_��lpWᐛ4�U���:!��	��g����k9����JLpդ��mw|-YB,E�sp_w��m���/�CR9�ﻺ�&Z��q�H����f3E���BR�����dMSI��Mf�h7ݩR;��ZS��w�%�z�J���48{�Uj��t�!�΄�|�D@���^�34��Mù��AY�3�qK7�N��9$�h]�#r�n�QAM�F�^����+�j��{���(���f�3���˃�r����������n���l�a!)B��mI��'U�v��z���������Ϻ�����E����n8s+���C��c��HX��E
����	�}�B� ��H�w�em���ԋ�j򰅥�`奲�?1����9F�%������g�0d*�mܡUH�U̢�M���,�5#�0�/��������@��F@j�3��&
.�Z�<{�= �����*z���S�"�)�7th�`F��|wġ������Qw�ڌbA?6�j�34�	�ѳ�E�5߲�J�l��y�`�/��gV@�9�e��Z��*�$�Ǜ���Y�?�j�vB���3cm�j0N��R��~��h�hoy�匽��3�&��[�\f�&;F�-"� ��5ph���k�j�[\�ua3o\���Z�Ó�D9���[!Q��g�'�M��=�����ө����2�Uo��<�Sj�ـc�k\:dW�o��]4q\f��}��Y�ؓ�-8���A�zN�ݐ�N,	�487|u�"Wn��� ߲hwQ�$�-	~z`�j����D�67�82�Т�����nI�_9�SC��L�*hb�h��Oȥf^��w�v�H�1�p�BA�i��-�W���n�Ö^
�~5���_¢U��@��G��&��;ޑ��M��N���2����6����{�o8_����}Y�/�Ϯɏ<�Ҍ4�d94�?�h+4������_�@}�dp5*�?a�~��0^���]	"��7���9h:l������A��z<�&״�~:-��!��?��4l�G�"y����}�De	4Q-�}�V��`���~��׏��/���bT}/��X��pd&ǡ;�0�����o�, M�Y���s1gL�=n���V��Lې��im�BPъ��ϕ�m��q\��`�@Ѝ���L�O:�=j
�T����7�#��FHb��1��&�Ϳ��|+����oʩ�rI"���kٕɱ�aL|��!���I'D{w�r��T��f!v|A'��c��m������
���6{x�K����h���Q�p�h�b����Ö�<��0>|�K�����G�[�)� �7+� ��W\�2f�J�h�T�HgA�.wp�+�3�&"^PB[�?sNOE<��P�y�%����r�6ڔ���`�^�S������z���mo�8�����ڋ��0)�'׼4-g�y�}��)+����1u+��VNK����K$�4� g����8����x�a��&��p�h��rW����A�����ߎ�'�C�+���~��@Ѳ�[�h����O��
p���i�AdVR�łO�d)cI�,�B[��n�	��~���-�v�H���L��Y�-�R���~%�f�(��;����N���Ҋ��A^+�Ŷڵn���P;���h��k�9GQ�غ��촢({ƨ�U��U&��|�������E�A$ ��j;�G	��	E�4So6������k6���Gذ�v��x���_"���ڙ�e��;޷ EQ�֪d 5��xDc��Q�V���X��y�ݶ�Dj���j\���Y ��o��a�C�N�m9��L���!�S0�K�(+kUc� @����͙�ks�X�{+�f�k��t��5�ƒ�R�B���dw����$�;U����
�����Ο���]v��g�ܳ~P[�������[��OB|�ߢ��|��v�N^u�D�i�����
�⁀	|Bl���]c�KKA3G���Y�W��������?$��I^�(pHG c�Cy��0�Z��)���Gy�rT��2�����e�/����,;hy�͝��8�?������q�Y9���9���+W��dN�,��1�r3W�h+��ޛ�'���}Ly����C�cO�1��-���$���#xJ�����b��?֜�v�(SRؐ\�j\���P~L��M��3�)�O���VR���Ĕ7��?��^���׸����6�4�4�x0�@�'7Sb��ʻ~�TF�I�*��0}b���_qe�ͪF�^����e�Iù�20m��U�/�4�K;D��Z�K$m�s��m�|llq�H٢�?Ek&U�� �m���^h�q��}�8�!(w���ex (�F��4��ϋ�9��S�L�j��������+�Z�%3}W���	p%�m��E<��7u��w,�+@��i�������v��\��[�UYm�k���n��t�5��Z������-8W�:�!32vOIǠm�ۈ����f�ⓛ<�}<��l,f��z���¬�%t��ÈC��\�IM"L>��Z��K�F�XQ�ƭ�=�8h8�k�a���p�t�����z09�M�'�����������*u��!1���`��j�v�K�x5l�7�?���H ���y�$����bl��&><E��0���dP@���m�1�I|dÛ�������t�1t���&V$%�����±������a/���-��NƒFq���\r��א��h 	�O��)�',���~�?�j�2�i��./�
kꙃvھl����Yh�q���3�cV_/f㫪��h`���#�	U����yK;����A[`R��P�p[��O��L�q��BF���|��j���P�N�q@8?"U>Q��aF����?��>�i���*˃�Q���8Z���NrȐ|�/�i"o>��ɜ��tx�Q^�������z�q-����r[|X��wqz7^1�$�1G UT���c,���u��%��+I��:A���♠�b�Ԗ}tUkߥ�iM��$s.�E�)��AJ*�oSr������X�aa%�nl�D�:��D20!�& #��*��S��k�_Z^�СS��
L�_뫆x���%  � &D��o���'H���8?�Zm��������we R���	��g�WX�]��q�f�(K=:"�]��Y����7�ɔ[d���T���=�g� �U_��d��Ș���aL�Ϫ�5��USI3O�o����ף{u;��Ӓo(���(V�a�CݳܗL+n��+O췟g�s��%Y��=lv�0$q)|��iv�-Wq�xw̯].��$;�ɦ��Cv�$�wM��A#B���<���r��5��蔦x�EÜ�������	�̄5�=l>���sR��%�����W\��(��w@��	~�lX�4=փ��ZY>�?��B����M�Щ��8K��Õ���B��ya]oV�A~�Wㄹ����Dې��X�C�%34�t͑e�A�����tUF�]6SN-�u<���{�F�<e�
��Gm�O�~1�h����8��}*��>!b�|�B9SkM6�ef6�C�����A�M{�`�/������t�>�o'����Aҙ?qT"]�����5j�����p�]�:d·s���8�əe[�}���пƶ��!���}ᏓL�a�0U�$x�)��7������aɸ�^-��`	�-/����n�k���D��\�Ns\��?ii�0UP�MK�ϖ��+b`g����m��od����$\�m�\X�l��/�˸��� �P�j�Pj�}ʷJ/�z3pWl*C�:7¡�I��Y;�����vsG���%���9\�Q��¿%�6'�Kg��ȣv�E^J0G��b��,Y��	(qƪf,���gy ��,�,��Q��Hm[�$1�ZX 3��` ���!Oi�|D�M/p?��c߮y*8d��u �R��A����!�co/�%q5d� ��6�㇒�)r��J\gy$5�>25�ײ���p�A�-��X���S���%�U�,�]�mq2�s̬f���2A�`	K�3�����Xk��>��J~ָ5����v8��j�I��ǩT���Qp��2rx�NM�.Kp���%��V ��V�c����zA<�CZ3�l�D[ؚ��g��b.������7�V������k 2��"�,k�]�'6����[!�m�����U�2��JZ���׀e��V3���p]�O �$6���]�4��藀�¿���d�GF���9���a�gw�^g�I��Xݦ~���X�yG�m#�z��X�9)$(�Zt�V����,��񰫉,�^�A�qԼ�Iq��*��4Bg�{�;:�N�D���!r�hnK�G+k�꽻�3mI���KbCe�!�A�@ch�ծe~	t�OS�,��].�&�a)�$ 0������sCcx�
u��!|P~N���I)8��'�z�k rS��X�=K�3rlrן�4M"E��ђA;jv��W�Gdk�	A�#�2���Ho���>�r�DCT�����PԻ0B�΢L�m������8厎Iڎ�'$.Ǟ���b����a�e�
P)�JUM�R��c��f�G��b�F}�#O�c ��U�v���ziH�[%5��Lu LA�W�u��{�>i��i�ݺ�lJEm�a��.�?ahڋ%U�$^��]�����C�k;aQI��-$����3G�dڜ��j��T:$����k�\��4Q �FB�=S0�$�ĹI��}'˫vW$ r	>�(g������f#[�ʿ�?�^0Sͱ�-��N-�A�n�q��g8�t(n{���'gU=f��k�M���� ��؛��o���:�H�=���e;�az7�U�*zIy��>m4xj(}�~�n�2� ��[ G+��! |e�モ֯��"l�	��}ut�G!W���H�tq
�������x�F����h!� ޷�smyy��xKUJ?i{���cc�/z��+W�V=0�5��K�U��7�v�ҷ6//1�0ڣ-S�R�8Ĭ��w�S��\�Z 5�ܥ�!D����il�V��2�K]B��&:��8��G���ρ]�i��{^;t��E�n7�S���S
3���{��Ʉ���ё�Vt�9���eY�XJv�G���"C�<Tn"�������ˠB� 1����#��4bП���R.w	�D�H�^�I=��j^=*��&�'�g�V�C)0K�ri֣A0�����u��
?�/��a�aGn'�^�%�{�ʯb{nm�[~��HD��p�+(}�+��W� c���-wv�v~sk ���6�[(Q���:q�S�RZ!��j��q|���`���z�I��lyb=}<?������p�ҫӌ��R38QWp���hT,���Q 辅v�r��[b0/�$�с�A�?��`�d�\��B<8�{H�� 
��9H �!]Lx���b����p�|�;��Qaj�&���-985��������Y� ?�X;m�*7)�y���&��?��犉'��ʽ�q�V����sі�?�﷫z����N,ŕ��@f�9CI���G�b=�>͒��\}f�P>q�scmq�Aj��A��w�E��ă��i�<ѽ�E����4�K� 1�Љ�de�^ZfM�5��w��tE�FA���甶#���"Ϲ�l� `G��cG.?��bw��A܇�0�C�s�y�-g#�QÞR���J�!�H㢾&���"u�ș�Ej�� ��'R(3�{@���e؊�Nd:oz�v �`��b�"�>�q�T��C���(�W2�;jc��ӕ��f���Mn>31,���G�5��2�RZY�l�'�b]IN5��Gϙ][�)����$)5��)P�;m�Y�;$��B\��1f%�IM��@�4t&�P�k���^;R@_��7p�X/��ǫ�N��!J��\;�p3V@�:�Om/��q����_�)k���E��p�v�x�k�@^�?�B�'�_���L]�(���?��L��q�]d���& I1��"j�t�j�$�����a3��&Ҙ���<�\�@�y���j48ց�Ĕ՛����޸����k��%2@�#)p��Kخ�פ�\Ϣ�	�����Z*ߠ���f���ړ�Xh_�ߎ�F0 ��B#�j/�wiKY���?��j�x�c⦱�m��FU�+��M��,L�(=���S���F||�`��p= S����σ���Ln�~>�}�ij�ɠO�"�_�[7p���I39�^_�:�@�� E3�`��;~@��Jws9��g}�]qX���+��2�/������R����^�F��J094=���x��o�@<�Ɩ3n�U��]G�6L�����J�J��/*;��C��)]#RAv&������B�DUT0�KE�~2����ђ�|un����ωգ�!�L�N��l�J�xۏXp%+O|��EnG�QJ8����۫_���%�+��+!�'�K����Т�n$X��W�T�=����O�g]:�O��i�%�Q���Ey�jR�
�6_'^����8{6x��)�Ȓǭ$ �/`�:��k�;���AVK��=�@��m,C+��7���pM���;f�n����!kF��_XT*QY�f��**�
��Hz�5�}�s]�;���By:cg����%�I$C��
� �X��R��ޝo������<�5s�
Mg�k��t��	��h��e�?z���7I��q0���*��NeR;�V���{bs)����V��.!?r����������*�q���eLm�CV����H.eP����/9��F
�n%]}�Y�h�8�`8(����% ����%,������#z�{5�7���&6�G����7�"�M0���g�ڎ��<9���tQ�91��vc]�G���0�;K�	�s�ޏz����0�J ���pr�G/�[�8��ķ�7�a1���svP)p��	��X�u�G�K&���a���|��c'>�k3����DU��T�7B5}ƃCm��.������s���Yn;U�l���*�E�Sf�C��4N!����"qOo�؋�9�G:,[?�y
V�5����^*뷽Ƚ#7����U�ؾX�I��4�^~Dif~��|P9~[�rƧ�����,��g�n��7�����d�M�Eu]�~k���ɒg�4K/l�
��.�O_�l���?4ۻl�ŷd���}��c	t0�3t�dS�j��1v.��UjT����:���K���87�cޕ����#�����zK���[���X���>
m�G?�4�S6ؒO= 9l�������b[�!DB	�$O
Ӯ�@���	�2�GV=s����˴{�H�!p�A~�ʂ` �*��j+N<�U���ʟ���=��aQyx��]-������k���e�v�������0^6i�B�9�׍j�t���
gg�BӘ�:���C/ߐ�]�8�t獕�Z���p�\�:٭���N�LH´5V4Eِw}R֟x�U0�\Ƥ�zD�'`3�A@����	a޲��ʞ-��_HP]�s��A��=��"�7Tؙ�?��m#��/�P����v���C�*[�1E�s�h�E�L�B���SoPd�&�Y,w��^�O�%"J��Tʷ�������/Ӹb�Z�9|`��}$��4��_�8��RV�w׋AZ�Pq�ϓOx��y��`�M�۲@E����s��L�kOg阾[�X���y��Fw�	ſkB���Z!i�Ϸ����^��"���(����YlK�KL��W:�6o|�|��܄)S���̢"{�_)c�P�̢�ՎeOo�S�{sSܿHM�(;�R��Cjɼӿ
�	6<�]�,8_Ѱ/C�!"E�e��\��S�;����Gv#F0�V���Ś�#c��ą����Ȟ�rtnmw0i�󨡤��a4���Q��(;T�n��: �h�]!�^?�L梽�]vaA"H�T�Jaޫ�{���h�-k��+�}��mJ���������)�Ų�F�:6��B��J^_=���h�a�U��SU�e��ڜگ��W�i��|�
Fj��Xm��4Dd7>~s������׮�![�.�i"L\� r��y��y���&E�kxr�������ypF�>�(�#�+�+ͦ��rJ�~s$p�R��-�F��Qo�"!�P�_5�1y�+je�f�֛�h�X�@�9��e�VdQ̖�~P>�c�f�ե�AvMy��÷ouP��aN�쾘z�9c��8h����%2Y�~�����t
��a�� ���C�����
�ş.����[Hq;��i���X��,��O=��L`!�����L���#��G��z|���$��ٲ�L�܇��:�9}���vZt�v�~|uD�i�B����nw)�=a��B����D�:zN�_�6�jӻ-v��*�y75S�i�[.�n^k#=v:�����2�G�NlT+�ݟּ��h�9rU&�G_���q����C��\�Fi�۔`�
j:Kɒ)�Ѥț<��Eļ_�I����$aB�;-�:D�N^}�@���R����"<u�*)�P���LlOk=e�C����|����% ���L�N1�]��<G��K�Y��S�Xwnw����[���eR��#�x0w�r 0����]ӕ���`�b]�b�8����gQ��;L�|H�߼c} u�w6׈;�y��g���s�~�@��;M�IM~��c�������p|�����
hy��x�eBЈ��N� �̧h���w�=c=1�̼_U=�L�Y��vP>z2ᣜ�L�tE�Cw\"AŚ<Z��ג�z����E����㟉����:�'��W9gƪ��s�<
�Z:��V�>m�R�Z�P���Z=�<<�O6Ζ��{��,Y���旃�y^	�'������V�
����Ő)����n�������F�`Fa�~)��/ET��ܳ�בk�/��b�4?L`FՇ�n�Y�2Ţ�|�*r�&"�+/E�y��v��.�˼
Cl����x�I� ��(@��c��8���)�~�=���j�ݣ����JbY0���Z�p'
xg>�R��>�aMn�|7� � Б��g
��}�|q]�HU_�u�{�s�����`D�*+,4Q&�iDU�`y�`;,�E��7��˕��~7�g�:O9���dZ�`oK��I��\W�P�(3�G�lo��EH����?j{�R���a9C��(*��3}f�*%�CP�m7�7����ԢP�����eZ?^/i�<��i�/]�����ޠ*׈vYbIX���� l2P[�=���)������Z��x#��1�-���Pw����b��՝o����7���=���Q��:vʒ<���D\�p=sN���
A��w�kf\~6��.�<`:I��0�(�؄��'���G���$m�u�����0A���G��	�p��cV-��჌�),��Sw�Г�W�������ԁ�_�t������P����P��������4�P,�g>0+O��O(S3((%F�V3ӕ��#��e�l{=�1*�g��7O�R���j���)�~��w6/�;J��n@+�(\+E��1q��0U�!��PLz�i��5.�B�10mc�b�6k�M��Z̰�&K�E�
0����	B'����<�Ie`�!E�-�ԙbi@����,x}:*�����$4h���~3�x�e��	r��^.�09�V��ή�Gw��*�VⷬYDj�ج`C�e߬�-Wƀ!xr��!HuPQ)Z�ʤt��pFC�{��Z㭿EF
Y~b��c˪(�	nh�=�g�D�����<��������-@�ο�R�:�7����p��j#���(d��I?[i�L7�\��sF\�����Jy��I[M���� <a{�v?k{�
�vQ)���L�"���Gh UU��j��$f�2��b�,��:�6!p�хa��&3|��4/K�,�M����k���"��psao;����L��Mjԥo*��